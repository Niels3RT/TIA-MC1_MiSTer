library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_g7 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_g7;

architecture rtl of rom_g7 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0000
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0008
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0010
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0018
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0020
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0028
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0038
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0048
         x"fb",  x"cc",  x"c6",  x"c6",  x"c6",  x"c6",  x"cc",  x"f8", -- 0050
         x"c3",  x"c0",  x"c0",  x"c0",  x"f8",  x"c0",  x"c0",  x"fe", -- 0058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0060
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0068
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0070
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0078
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0080
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0088
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0090
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0098
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00D0
         x"01",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe", -- 00D8
         x"c0",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf", -- 00E0
         x"ff",  x"ff",  x"ff",  x"cf",  x"f7",  x"07",  x"1f",  x"0c", -- 00E8
         x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"01", -- 00F0
         x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"c0", -- 00F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0100
         x"c8",  x"e1",  x"33",  x"f7",  x"ef",  x"ff",  x"ff",  x"ff", -- 0108
         x"f8",  x"ff",  x"fe",  x"fe",  x"fe",  x"ff",  x"ff",  x"ff", -- 0110
         x"7f",  x"7f",  x"bf",  x"cf",  x"e3",  x"e0",  x"e0",  x"f0", -- 0118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"f8",  x"f0",  x"c0", -- 0130
         x"ff",  x"ff",  x"7f",  x"7f",  x"3f",  x"1f",  x"0f",  x"03", -- 0138
         x"44",  x"44",  x"44",  x"44",  x"44",  x"44",  x"44",  x"44", -- 0140
         x"44",  x"44",  x"44",  x"44",  x"00",  x"00",  x"00",  x"00", -- 0148
         x"ff",  x"ff",  x"7f",  x"7f",  x"3f",  x"1f",  x"0f",  x"03", -- 0150
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"f8",  x"f0",  x"c0", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0160
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"7f",  x"3f",  x"1f",  x"0f",  x"07",  x"03",  x"01",  x"00", -- 0170
         x"7e",  x"02",  x"02",  x"00",  x"e7",  x"20",  x"20",  x"00", -- 0178
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0180
         x"1c",  x"08",  x"1c",  x"3c",  x"9e",  x"0c",  x"14",  x"42", -- 0188
         x"01",  x"02",  x"04",  x"08",  x"10",  x"20",  x"40",  x"80", -- 0190
         x"80",  x"40",  x"20",  x"10",  x"08",  x"04",  x"02",  x"01", -- 0198
         x"80",  x"40",  x"20",  x"10",  x"08",  x"04",  x"02",  x"01", -- 01A0
         x"01",  x"02",  x"04",  x"08",  x"10",  x"20",  x"40",  x"80", -- 01A8
         x"fe",  x"fc",  x"f8",  x"f0",  x"e0",  x"c0",  x"80",  x"00", -- 01B0
         x"00",  x"00",  x"00",  x"00",  x"18",  x"18",  x"3c",  x"7e", -- 01B8
         x"00",  x"77",  x"77",  x"77",  x"77",  x"77",  x"77",  x"00", -- 01C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D0
         x"00",  x"03",  x"0f",  x"1f",  x"3f",  x"ff",  x"ff",  x"ff", -- 01D8
         x"10",  x"00",  x"00",  x"02",  x"07",  x"07",  x"0f",  x"9f", -- 01E0
         x"08",  x"c0",  x"c4",  x"ee",  x"ff",  x"ff",  x"ff",  x"ff", -- 01E8
         x"00",  x"00",  x"02",  x"07",  x"27",  x"7f",  x"7f",  x"7f", -- 01F0
         x"00",  x"80",  x"c0",  x"e8",  x"ec",  x"fc",  x"fc",  x"fe", -- 01F8
         x"ff",  x"fc",  x"f8",  x"f0",  x"e0",  x"e0",  x"c0",  x"80", -- 0200
         x"00",  x"00",  x"00",  x"04",  x"3e",  x"7e",  x"ff",  x"ff", -- 0208
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0210
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0218
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0220
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0228
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0230
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0238
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0240
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0248
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0250
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0258
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0260
         x"fe",  x"fc",  x"f8",  x"f0",  x"e0",  x"c0",  x"c0",  x"87", -- 0268
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0270
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0278
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0280
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0288
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0290
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0298
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0300
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0308
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0310
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0318
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0320
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"0f", -- 0328
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"e0", -- 0330
         x"0f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0338
         x"e0",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0340
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0348
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0350
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0358
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"0f",  x"ff",  x"3c", -- 0360
         x"e7",  x"f7",  x"ff",  x"ff",  x"ff",  x"fe",  x"ff",  x"f8", -- 0368
         x"0f",  x"e3",  x"ff",  x"ff",  x"ff",  x"f1",  x"ff",  x"e1", -- 0370
         x"80",  x"c3",  x"ff",  x"ff",  x"ff",  x"c4",  x"ff",  x"c3", -- 0378
         x"9f",  x"ff",  x"ef",  x"ff",  x"ff",  x"ff",  x"f1",  x"e0", -- 0380
         x"f1",  x"ff",  x"c3",  x"ff",  x"ff",  x"ff",  x"cf",  x"e7", -- 0388
         x"c3",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"e3",  x"07", -- 0390
         x"c3",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c3",  x"80", -- 0398
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"ff",  x"7f", -- 03A0
         x"83",  x"c7",  x"ff",  x"ff",  x"ff",  x"c4",  x"ff",  x"c4", -- 03A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03B0
         x"83",  x"c7",  x"ff",  x"ff",  x"ff",  x"c7",  x"ff",  x"c7", -- 03B8
         x"0f",  x"ff",  x"f1",  x"ff",  x"ff",  x"ff",  x"e1",  x"07", -- 03C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"e3",  x"07", -- 03D0
         x"c7",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c3",  x"80", -- 03D8
         x"1f",  x"07",  x"ff",  x"ff",  x"ff",  x"f8",  x"ff",  x"ff", -- 03E0
         x"f8",  x"e0",  x"ff",  x"ff",  x"ff",  x"1c",  x"ff",  x"3b", -- 03E8
         x"c1",  x"e3",  x"ff",  x"ff",  x"ff",  x"e3",  x"ff",  x"e3", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F8
         x"ff",  x"ff",  x"00",  x"ff",  x"ff",  x"ff",  x"0f",  x"1f", -- 0400
         x"3c",  x"ff",  x"3e",  x"ff",  x"ff",  x"ff",  x"e0",  x"f8", -- 0408
         x"c3",  x"ff",  x"03",  x"ff",  x"ff",  x"ff",  x"e3",  x"c1", -- 0410
         x"c1",  x"ff",  x"c6",  x"ff",  x"ff",  x"ff",  x"c7",  x"f3", -- 0418
         x"1f",  x"07",  x"ff",  x"ff",  x"ff",  x"fc",  x"ff",  x"fc", -- 0420
         x"f8",  x"e0",  x"ff",  x"ff",  x"ff",  x"1f",  x"ff",  x"3f", -- 0428
         x"e0",  x"f1",  x"ff",  x"ff",  x"ff",  x"e3",  x"ff",  x"e1", -- 0430
         x"83",  x"c7",  x"ff",  x"ff",  x"ff",  x"c4",  x"ff",  x"c3", -- 0438
         x"fc",  x"ff",  x"f8",  x"ff",  x"ff",  x"ff",  x"07",  x"1f", -- 0440
         x"3f",  x"ff",  x"3f",  x"ff",  x"ff",  x"ff",  x"e0",  x"f8", -- 0448
         x"c5",  x"ff",  x"07",  x"ff",  x"ff",  x"ff",  x"f0",  x"e0", -- 0450
         x"c3",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c7",  x"f3", -- 0458
         x"ff",  x"ff",  x"7f",  x"3f",  x"07",  x"03",  x"19",  x"3c", -- 0460
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0468
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0470
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0478
         x"01",  x"01",  x"00",  x"06",  x"fe",  x"f8",  x"00",  x"00", -- 0480
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0488
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"00", -- 0490
         x"a6",  x"78",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0498
         x"01",  x"ab",  x"bd",  x"60",  x"e0",  x"80",  x"00",  x"00", -- 04A0
         x"00",  x"80",  x"80",  x"60",  x"7f",  x"1f",  x"00",  x"00", -- 04A8
         x"00",  x"00",  x"00",  x"80",  x"80",  x"80",  x"80",  x"00", -- 04B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 04B8
         x"b4",  x"dd",  x"eb",  x"07",  x"03",  x"00",  x"00",  x"00", -- 04C0
         x"92",  x"76",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 04C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"ff", -- 04D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fd",  x"ff", -- 04D8
         x"1f",  x"5f",  x"1f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 04E0
         x"f1",  x"f3",  x"f1",  x"fd",  x"ff",  x"ff",  x"ff",  x"ff", -- 04E8
         x"01",  x"00",  x"40",  x"04",  x"00",  x"10",  x"02",  x"00", -- 04F0
         x"80",  x"c0",  x"c0",  x"60",  x"04",  x"04",  x"06",  x"00", -- 04F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0500
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0508
         x"f8",  x"e3",  x"ef",  x"ef",  x"8f",  x"bf",  x"3f",  x"7f", -- 0510
         x"ff",  x"ff",  x"ff",  x"ff",  x"e1",  x"c8",  x"9c",  x"3e", -- 0518
         x"01",  x"07",  x"1f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 0520
         x"00",  x"00",  x"00",  x"00",  x"01",  x"07",  x"1f",  x"7f", -- 0528
         x"01",  x"00",  x"10",  x"30",  x"30",  x"10",  x"00",  x"00", -- 0530
         x"c7",  x"93",  x"bf",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0538
         x"ff",  x"75",  x"a5",  x"14",  x"02",  x"00",  x"00",  x"00", -- 0540
         x"00",  x"8a",  x"5a",  x"eb",  x"fd",  x"ff",  x"ff",  x"ff", -- 0548
         x"ff",  x"75",  x"a5",  x"14",  x"02",  x"00",  x"00",  x"b9", -- 0550
         x"01",  x"05",  x"05",  x"0f",  x"0a",  x"00",  x"01",  x"03", -- 0558
         x"78",  x"34",  x"14",  x"18",  x"34",  x"64",  x"64",  x"74", -- 0560
         x"00",  x"02",  x"03",  x"07",  x"07",  x"05",  x"01",  x"00", -- 0568
         x"78",  x"60",  x"2c",  x"3e",  x"1a",  x"32",  x"52",  x"50", -- 0570
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0578
         x"00",  x"00",  x"00",  x"00",  x"80",  x"e0",  x"f8",  x"fe", -- 0580
         x"80",  x"e0",  x"f8",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff", -- 0588
         x"ff",  x"ff",  x"ff",  x"ff",  x"e3",  x"c3",  x"80",  x"00", -- 0590
         x"00",  x"80",  x"c0",  x"e0",  x"f0",  x"f8",  x"fc",  x"fe", -- 0598
         x"00",  x"80",  x"e0",  x"f8",  x"fe",  x"ff",  x"ff",  x"ff", -- 05A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"83",  x"c7",  x"ff", -- 05A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 05B0
         x"ff",  x"7f",  x"3f",  x"9f",  x"df",  x"c3",  x"f0",  x"fc", -- 05B8
         x"ff",  x"ff",  x"ff",  x"fc",  x"f9",  x"83",  x"bf",  x"7f", -- 05C0
         x"fc",  x"fe",  x"fe",  x"e6",  x"c0",  x"e0",  x"c0",  x"00", -- 05C8
         x"ff",  x"8f",  x"2f",  x"e3",  x"f1",  x"fd",  x"fc",  x"fe", -- 05D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 05D8
         x"cf",  x"9f",  x"9f",  x"3f",  x"3f",  x"9e",  x"cd",  x"e3", -- 05E0
         x"c3",  x"9d",  x"3e",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 05E8
         x"e3",  x"ca",  x"dc",  x"9f",  x"9f",  x"3f",  x"7f",  x"7f", -- 05F0
         x"00",  x"1c",  x"3e",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 05F8
         x"00",  x"03",  x"0f",  x"3f",  x"ff",  x"ff",  x"ff",  x"ff", -- 0600
         x"00",  x"01",  x"03",  x"07",  x"0f",  x"1f",  x"3f",  x"7f", -- 0608
         x"ff",  x"ff",  x"ff",  x"ff",  x"ef",  x"c3",  x"98",  x"3c", -- 0610
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0618
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0620
         x"e3",  x"c9",  x"9c",  x"3f",  x"ff",  x"ff",  x"ff",  x"ff", -- 0628
         x"fc",  x"fe",  x"f2",  x"e0",  x"e0",  x"e0",  x"80",  x"00", -- 0630
         x"00",  x"18",  x"3c",  x"fe",  x"fe",  x"fe",  x"fc",  x"f8", -- 0638
         x"f9",  x"f0",  x"f6",  x"e7",  x"8f",  x"3f",  x"7f",  x"3f", -- 0640
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0648
         x"3f",  x"1f",  x"1f",  x"0f",  x"61",  x"7c",  x"7f",  x"ff", -- 0650
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f", -- 0658
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0660
         x"ff",  x"ff",  x"ff",  x"77",  x"23",  x"03",  x"03",  x"00", -- 0668
         x"ff",  x"ff",  x"ff",  x"fe",  x"fc",  x"f8",  x"60",  x"00", -- 0670
         x"00",  x"00",  x"02",  x"06",  x"1f",  x"1f",  x"3f",  x"1f", -- 0678
         x"ff",  x"ff",  x"ff",  x"1f",  x"0f",  x"07",  x"00",  x"00", -- 0680
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0688
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0690
         x"c7",  x"9f",  x"3e",  x"7e",  x"3e",  x"bf",  x"9f",  x"cf", -- 0698
         x"00",  x"00",  x"00",  x"00",  x"00",  x"1c",  x"3f",  x"7e", -- 06A0
         x"80",  x"e0",  x"f8",  x"c0",  x"f0",  x"fc",  x"fe",  x"ff", -- 06A8
         x"00",  x"18",  x"3c",  x"3e",  x"ff",  x"ff",  x"ff",  x"ff", -- 06B0
         x"0f",  x"03",  x"03",  x"01",  x"00",  x"00",  x"00",  x"00", -- 06B8
         x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe", -- 06C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 06C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 06E0
         x"f8",  x"70",  x"90",  x"08",  x"00",  x"00",  x"80",  x"e0", -- 06E8
         x"83",  x"8f",  x"7f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 06F0
         x"f0",  x"f8",  x"fc",  x"de",  x"bf",  x"9f",  x"c7",  x"ff", -- 06F8
         x"00",  x"00",  x"09",  x"1f",  x"03",  x"07",  x"0f",  x"0f", -- 0700
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0708
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0710
         x"1f",  x"bf",  x"bf",  x"bf",  x"bf",  x"ff",  x"ff",  x"ff", -- 0718
         x"00",  x"88",  x"cd",  x"dd",  x"dd",  x"fd",  x"ff",  x"ff", -- 0720
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0728
         x"1f",  x"07",  x"f3",  x"f3",  x"fb",  x"f9",  x"fc",  x"ff", -- 0730
         x"e7",  x"f3",  x"fb",  x"fd",  x"fd",  x"f9",  x"f3",  x"07", -- 0738
         x"fe",  x"fe",  x"fe",  x"fd",  x"fd",  x"f3",  x"cf",  x"1f", -- 0740
         x"fe",  x"fe",  x"fe",  x"ed",  x"d3",  x"ef",  x"cf",  x"3f", -- 0748
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0750
         x"7f",  x"3f",  x"b7",  x"83",  x"cb",  x"fb",  x"f8",  x"fe", -- 0758
         x"e7",  x"cf",  x"9f",  x"df",  x"df",  x"cf",  x"e3",  x"f8", -- 0760
         x"ff",  x"ff",  x"ff",  x"ff",  x"ec",  x"c0",  x"c0",  x"00", -- 0768
         x"ff",  x"ff",  x"7f",  x"3f",  x"07",  x"03",  x"01",  x"00", -- 0770
         x"f8",  x"fc",  x"fe",  x"fe",  x"ee",  x"c4",  x"c0",  x"00", -- 0778
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0780
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0788
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0790
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0800
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0808
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0810
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0818
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0820
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0828
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80", -- 0830
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80", -- 0838
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 0840
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"ff", -- 0848
         x"fb",  x"cc",  x"c6",  x"c6",  x"c6",  x"c6",  x"cc",  x"f8", -- 0850
         x"c3",  x"c0",  x"c0",  x"c0",  x"f8",  x"c0",  x"c0",  x"fe", -- 0858
         x"80",  x"80",  x"80",  x"88",  x"80",  x"80",  x"80",  x"ff", -- 0860
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0868
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0870
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0878
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0880
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0888
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0890
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0898
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08C8
         x"fe",  x"f9",  x"e3",  x"83",  x"07",  x"3f",  x"7f",  x"ff", -- 08D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f", -- 08E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 08F8
         x"fa",  x"f7",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0900
         x"ff",  x"ff",  x"df",  x"cf",  x"ff",  x"3f",  x"1f",  x"3f", -- 0908
         x"f8",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"ff", -- 0910
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"ff",  x"fc", -- 0918
         x"ff",  x"ff",  x"fe",  x"fe",  x"ff",  x"ff",  x"f7",  x"c0", -- 0920
         x"ff",  x"ff",  x"7f",  x"7f",  x"ff",  x"ff",  x"ef",  x"03", -- 0928
         x"ff",  x"ff",  x"fe",  x"fe",  x"ff",  x"ff",  x"f7",  x"c0", -- 0930
         x"ff",  x"ff",  x"7f",  x"7f",  x"ff",  x"ff",  x"ef",  x"03", -- 0938
         x"7e",  x"7e",  x"7e",  x"44",  x"e7",  x"e7",  x"e7",  x"44", -- 0940
         x"7e",  x"7e",  x"7e",  x"44",  x"e7",  x"ef",  x"e7",  x"44", -- 0948
         x"ff",  x"ff",  x"7f",  x"7f",  x"3f",  x"1f",  x"0f",  x"03", -- 0950
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"f8",  x"f0",  x"c0", -- 0958
         x"00",  x"00",  x"01",  x"00",  x"03",  x"07",  x"07",  x"00", -- 0960
         x"00",  x"00",  x"80",  x"00",  x"c0",  x"e0",  x"e0",  x"00", -- 0968
         x"7f",  x"3f",  x"1f",  x"0f",  x"07",  x"03",  x"01",  x"00", -- 0970
         x"7e",  x"02",  x"02",  x"00",  x"e7",  x"20",  x"20",  x"00", -- 0978
         x"7e",  x"7e",  x"7e",  x"00",  x"ef",  x"ef",  x"ef",  x"1c", -- 0980
         x"7e",  x"7e",  x"7e",  x"3c",  x"ff",  x"ef",  x"f7",  x"42", -- 0988
         x"7f",  x"7e",  x"7e",  x"08",  x"f7",  x"e7",  x"e7",  x"80", -- 0990
         x"fe",  x"7e",  x"7e",  x"10",  x"ef",  x"e7",  x"e7",  x"01", -- 0998
         x"fe",  x"7e",  x"7f",  x"17",  x"ef",  x"f7",  x"e7",  x"01", -- 09A0
         x"7f",  x"7e",  x"f4",  x"ef",  x"f7",  x"ef",  x"e7",  x"80", -- 09A8
         x"fe",  x"fc",  x"f8",  x"f0",  x"e0",  x"c0",  x"80",  x"00", -- 09B0
         x"e7",  x"e7",  x"e7",  x"00",  x"ff",  x"ff",  x"3c",  x"ff", -- 09B8
         x"00",  x"77",  x"77",  x"77",  x"77",  x"77",  x"77",  x"00", -- 09C0
         x"00",  x"7c",  x"7c",  x"00",  x"00",  x"c7",  x"c7",  x"00", -- 09C8
         x"77",  x"3f",  x"7f",  x"7f",  x"4b",  x"c0",  x"00",  x"00", -- 09D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 09D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 09E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 09E8
         x"00",  x"00",  x"02",  x"07",  x"27",  x"7f",  x"7f",  x"7f", -- 09F0
         x"00",  x"80",  x"c0",  x"e8",  x"ec",  x"fc",  x"fc",  x"fe", -- 09F8
         x"ff",  x"fc",  x"f8",  x"f0",  x"e0",  x"e0",  x"c0",  x"80", -- 0A00
         x"00",  x"04",  x"3f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"01",  x"07",  x"00", -- 0A68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0AF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"0f", -- 0B28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"e0", -- 0B30
         x"0f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B38
         x"e0",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"3c", -- 0B60
         x"e7",  x"ff",  x"ff",  x"ff",  x"fc",  x"ff",  x"ff",  x"f8", -- 0B68
         x"0f",  x"ff",  x"ff",  x"ff",  x"f1",  x"ff",  x"ff",  x"e1", -- 0B70
         x"80",  x"ff",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"c3", -- 0B78
         x"9f",  x"ff",  x"ff",  x"e7",  x"ff",  x"ff",  x"ff",  x"e0", -- 0B80
         x"f1",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"e7", -- 0B88
         x"c3",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"07", -- 0B90
         x"c3",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"80", -- 0B98
         x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"ff",  x"ff",  x"7f", -- 0BA0
         x"83",  x"ff",  x"ff",  x"ff",  x"c6",  x"ff",  x"ff",  x"c4", -- 0BA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BB0
         x"83",  x"ff",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"c7", -- 0BB8
         x"0f",  x"ff",  x"ff",  x"f1",  x"ff",  x"ff",  x"ff",  x"07", -- 0BC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"07", -- 0BD0
         x"c7",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"80", -- 0BD8
         x"1f",  x"ff",  x"ff",  x"ff",  x"f9",  x"ff",  x"ff",  x"ff", -- 0BE0
         x"f8",  x"ff",  x"ff",  x"ff",  x"8f",  x"ff",  x"ff",  x"3b", -- 0BE8
         x"c1",  x"ff",  x"ff",  x"ff",  x"e3",  x"ff",  x"ff",  x"e3", -- 0BF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BF8
         x"ff",  x"ff",  x"ff",  x"f1",  x"ff",  x"ff",  x"ff",  x"1f", -- 0C00
         x"3c",  x"ff",  x"ff",  x"bf",  x"ff",  x"ff",  x"ff",  x"f8", -- 0C08
         x"c3",  x"ff",  x"ff",  x"e3",  x"ff",  x"ff",  x"ff",  x"c1", -- 0C10
         x"c1",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"f3", -- 0C18
         x"1f",  x"ff",  x"ff",  x"ff",  x"fd",  x"ff",  x"ff",  x"fc", -- 0C20
         x"f8",  x"ff",  x"ff",  x"ff",  x"8f",  x"ff",  x"ff",  x"3f", -- 0C28
         x"e0",  x"ff",  x"ff",  x"ff",  x"e3",  x"ff",  x"ff",  x"e1", -- 0C30
         x"83",  x"ff",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"c3", -- 0C38
         x"fc",  x"ff",  x"ff",  x"f1",  x"ff",  x"ff",  x"ff",  x"1f", -- 0C40
         x"3f",  x"ff",  x"ff",  x"bf",  x"ff",  x"ff",  x"ff",  x"f8", -- 0C48
         x"c5",  x"ff",  x"ff",  x"e3",  x"ff",  x"ff",  x"ff",  x"e0", -- 0C50
         x"c3",  x"ff",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"f3", -- 0C58
         x"00",  x"00",  x"80",  x"c0",  x"f8",  x"fc",  x"fe",  x"ff", -- 0C60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C78
         x"01",  x"01",  x"01",  x"07",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff", -- 0C90
         x"59",  x"84",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C98
         x"fe",  x"54",  x"42",  x"80",  x"00",  x"00",  x"00",  x"00", -- 0CA0
         x"00",  x"80",  x"80",  x"e0",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CA8
         x"00",  x"00",  x"00",  x"80",  x"80",  x"80",  x"80",  x"00", -- 0CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 0CB8
         x"4b",  x"22",  x"14",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CC0
         x"6d",  x"09",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CC8
         x"ff",  x"7f",  x"1f",  x"0f",  x"cf",  x"0f",  x"07",  x"07", -- 0CD0
         x"ff",  x"fc",  x"f0",  x"e1",  x"e7",  x"e0",  x"c0",  x"c0", -- 0CD8
         x"23",  x"63",  x"e3",  x"83",  x"03",  x"07",  x"0f",  x"1f", -- 0CE0
         x"88",  x"8a",  x"8e",  x"82",  x"80",  x"c0",  x"e0",  x"f8", -- 0CE8
         x"01",  x"00",  x"40",  x"04",  x"00",  x"10",  x"02",  x"00", -- 0CF0
         x"e0",  x"f0",  x"f0",  x"e0",  x"4e",  x"0f",  x"06",  x"ff", -- 0CF8
         x"00",  x"80",  x"c1",  x"c1",  x"c3",  x"e3",  x"e3",  x"f7", -- 0D00
         x"01",  x"07",  x"01",  x"03",  x"07",  x"03",  x"07",  x"0f", -- 0D08
         x"07",  x"1c",  x"10",  x"10",  x"70",  x"40",  x"c0",  x"80", -- 0D10
         x"00",  x"00",  x"00",  x"00",  x"1e",  x"37",  x"63",  x"c1", -- 0D18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D28
         x"03",  x"03",  x"79",  x"fd",  x"fc",  x"78",  x"00",  x"ff", -- 0D30
         x"b8",  x"ec",  x"c0",  x"80",  x"00",  x"00",  x"80",  x"80", -- 0D38
         x"00",  x"8a",  x"5a",  x"eb",  x"fd",  x"ff",  x"ff",  x"ff", -- 0D40
         x"ff",  x"75",  x"a5",  x"14",  x"02",  x"00",  x"00",  x"00", -- 0D48
         x"00",  x"8a",  x"5a",  x"eb",  x"fd",  x"ff",  x"ff",  x"46", -- 0D50
         x"2f",  x"6f",  x"7f",  x"df",  x"df",  x"4f",  x"6f",  x"0f", -- 0D58
         x"78",  x"34",  x"14",  x"18",  x"34",  x"64",  x"64",  x"74", -- 0D60
         x"5f",  x"5f",  x"3f",  x"3f",  x"5f",  x"0f",  x"af",  x"af", -- 0D68
         x"78",  x"60",  x"2c",  x"3e",  x"1a",  x"32",  x"52",  x"50", -- 0D70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D78
         x"00",  x"03",  x"07",  x"03",  x"81",  x"e1",  x"f8",  x"fe", -- 0D80
         x"80",  x"e0",  x"f8",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D88
         x"00",  x"00",  x"00",  x"00",  x"1c",  x"3c",  x"67",  x"c3", -- 0D90
         x"00",  x"80",  x"c0",  x"e0",  x"f0",  x"f8",  x"fc",  x"fe", -- 0D98
         x"07",  x"81",  x"e1",  x"f8",  x"fe",  x"ff",  x"ff",  x"ff", -- 0DA0
         x"ff",  x"ff",  x"ff",  x"7f",  x"3f",  x"9f",  x"df",  x"ff", -- 0DA8
         x"07",  x"8f",  x"9f",  x"df",  x"df",  x"df",  x"df",  x"ff", -- 0DB0
         x"00",  x"80",  x"c0",  x"e0",  x"e0",  x"fc",  x"ff",  x"ff", -- 0DB8
         x"00",  x"00",  x"00",  x"03",  x"07",  x"7f",  x"7f",  x"ff", -- 0DC0
         x"03",  x"01",  x"01",  x"19",  x"26",  x"10",  x"20",  x"c0", -- 0DC8
         x"ff",  x"ff",  x"df",  x"1f",  x"0f",  x"03",  x"03",  x"01", -- 0DD0
         x"00",  x"8c",  x"d8",  x"dc",  x"fe",  x"fc",  x"fe",  x"ff", -- 0DD8
         x"f0",  x"e0",  x"e0",  x"c0",  x"c0",  x"e1",  x"f3",  x"ff", -- 0DE0
         x"ff",  x"e3",  x"c1",  x"80",  x"00",  x"00",  x"00",  x"00", -- 0DE8
         x"ff",  x"f7",  x"e3",  x"e0",  x"e0",  x"c0",  x"80",  x"80", -- 0DF0
         x"3c",  x"62",  x"c1",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E08
         x"00",  x"00",  x"00",  x"00",  x"10",  x"3c",  x"7f",  x"ff", -- 0E10
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"f8",  x"e0",  x"80", -- 0E18
         x"fe",  x"f8",  x"e0",  x"80",  x"00",  x"00",  x"00",  x"00", -- 0E20
         x"1c",  x"36",  x"63",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 0E28
         x"02",  x"01",  x"0d",  x"16",  x"10",  x"18",  x"60",  x"80", -- 0E30
         x"38",  x"64",  x"c2",  x"01",  x"01",  x"01",  x"02",  x"04", -- 0E38
         x"ff",  x"ff",  x"f9",  x"f8",  x"f0",  x"c0",  x"80",  x"c0", -- 0E40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E58
         x"00",  x"00",  x"80",  x"e0",  x"00",  x"c0",  x"f0",  x"c0", -- 0E60
         x"00",  x"00",  x"00",  x"88",  x"dc",  x"6c",  x"0c",  x"07", -- 0E68
         x"00",  x"00",  x"00",  x"01",  x"02",  x"04",  x"9c",  x"e0", -- 0E70
         x"00",  x"07",  x"1d",  x"39",  x"60",  x"60",  x"c0",  x"e0", -- 0E78
         x"00",  x"00",  x"00",  x"e0",  x"30",  x"18",  x"0f",  x"03", -- 0E80
         x"01",  x"0f",  x"03",  x"07",  x"1f",  x"07",  x"0f",  x"3f", -- 0E88
         x"00",  x"01",  x"0f",  x"07",  x"01",  x"1f",  x"03",  x"00", -- 0E90
         x"38",  x"60",  x"c0",  x"80",  x"c0",  x"40",  x"60",  x"30", -- 0E98
         x"e0",  x"f0",  x"c0",  x"fc",  x"f0",  x"fc",  x"ff",  x"fe", -- 0EA0
         x"80",  x"e0",  x"f8",  x"c0",  x"f0",  x"fc",  x"fe",  x"ff", -- 0EA8
         x"3c",  x"66",  x"43",  x"c1",  x"00",  x"00",  x"00",  x"00", -- 0EB0
         x"70",  x"1c",  x"0c",  x"0e",  x"03",  x"01",  x"01",  x"00", -- 0EB8
         x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe", -- 0EC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EC8
         x"00",  x"80",  x"e0",  x"c0",  x"f8",  x"e0",  x"e0",  x"80", -- 0ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EE0
         x"07",  x"83",  x"41",  x"c3",  x"e3",  x"e3",  x"f1",  x"fc", -- 0EE8
         x"7f",  x"7c",  x"f0",  x"e0",  x"c0",  x"c0",  x"80",  x"80", -- 0EF0
         x"ff",  x"3f",  x"0f",  x"27",  x"43",  x"63",  x"39",  x"01", -- 0EF8
         x"00",  x"00",  x"09",  x"1f",  x"03",  x"07",  x"0f",  x"0f", -- 0F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0F10
         x"1f",  x"bf",  x"bf",  x"bf",  x"bf",  x"ff",  x"ff",  x"ff", -- 0F18
         x"00",  x"88",  x"cd",  x"dd",  x"dd",  x"fd",  x"ff",  x"ff", -- 0F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0F28
         x"e0",  x"f8",  x"0c",  x"0c",  x"04",  x"06",  x"03",  x"00", -- 0F30
         x"18",  x"0c",  x"04",  x"02",  x"02",  x"06",  x"0c",  x"f8", -- 0F38
         x"01",  x"01",  x"01",  x"02",  x"02",  x"0c",  x"30",  x"e0", -- 0F40
         x"01",  x"01",  x"01",  x"12",  x"2c",  x"10",  x"30",  x"c0", -- 0F48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0F50
         x"80",  x"c0",  x"48",  x"7c",  x"34",  x"04",  x"07",  x"01", -- 0F58
         x"18",  x"30",  x"60",  x"20",  x"20",  x"30",  x"1c",  x"07", -- 0F60
         x"00",  x"00",  x"00",  x"00",  x"13",  x"2c",  x"20",  x"c0", -- 0F68
         x"00",  x"00",  x"80",  x"c0",  x"78",  x"0c",  x"06",  x"03", -- 0F70
         x"04",  x"02",  x"01",  x"01",  x"11",  x"3a",  x"2c",  x"c0", -- 0F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0F88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1000
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1008
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1010
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1018
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1020
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1028
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80", -- 1030
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80", -- 1038
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 1040
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"ff", -- 1048
         x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1050
         x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1058
         x"80",  x"80",  x"80",  x"88",  x"80",  x"80",  x"80",  x"ff", -- 1060
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1068
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1070
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1078
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1080
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1088
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1090
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1098
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f", -- 10E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10F8
         x"fa",  x"f7",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1100
         x"bf",  x"df",  x"ef",  x"7f",  x"7f",  x"ff",  x"ff",  x"ff", -- 1108
         x"f8",  x"f0",  x"f9",  x"fd",  x"fd",  x"ff",  x"ff",  x"ff", -- 1110
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7e",  x"5f",  x"bc", -- 1118
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1120
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1128
         x"00",  x"00",  x"01",  x"01",  x"03",  x"07",  x"0f",  x"3f", -- 1130
         x"00",  x"00",  x"80",  x"80",  x"c0",  x"e0",  x"f0",  x"fc", -- 1138
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1140
         x"ff",  x"ff",  x"ff",  x"ff",  x"bb",  x"11",  x"bb",  x"bb", -- 1148
         x"ff",  x"ff",  x"7f",  x"7f",  x"3f",  x"1f",  x"0f",  x"03", -- 1150
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"f8",  x"f0",  x"c0", -- 1158
         x"00",  x"00",  x"01",  x"01",  x"03",  x"07",  x"0f",  x"3f", -- 1160
         x"00",  x"00",  x"80",  x"80",  x"c0",  x"e0",  x"f0",  x"fc", -- 1168
         x"80",  x"80",  x"80",  x"f0",  x"18",  x"18",  x"18",  x"ff", -- 1170
         x"ff",  x"83",  x"83",  x"ff",  x"ff",  x"38",  x"38",  x"ff", -- 1178
         x"f7",  x"f7",  x"f7",  x"e3",  x"f7",  x"f7",  x"f7",  x"e3", -- 1180
         x"ff",  x"f7",  x"e3",  x"c3",  x"61",  x"f3",  x"eb",  x"bd", -- 1188
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1190
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1198
         x"c3",  x"f1",  x"f0",  x"f8",  x"dc",  x"ef",  x"ff",  x"ff", -- 11A0
         x"c3",  x"8f",  x"0f",  x"1f",  x"3b",  x"f7",  x"ff",  x"ff", -- 11A8
         x"01",  x"01",  x"01",  x"0f",  x"08",  x"08",  x"08",  x"ff", -- 11B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"e7",  x"e7",  x"c3",  x"81", -- 11B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 11C0
         x"81",  x"fd",  x"fd",  x"ff",  x"18",  x"df",  x"df",  x"ff", -- 11C8
         x"77",  x"35",  x"50",  x"00",  x"34",  x"3f",  x"ff",  x"ff", -- 11D0
         x"ff",  x"fc",  x"f0",  x"e0",  x"c0",  x"00",  x"00",  x"00", -- 11D8
         x"ef",  x"ff",  x"ff",  x"fd",  x"f8",  x"f8",  x"f0",  x"60", -- 11E0
         x"f7",  x"3f",  x"3b",  x"11",  x"00",  x"00",  x"00",  x"00", -- 11E8
         x"ff",  x"ff",  x"fd",  x"f8",  x"d8",  x"80",  x"80",  x"80", -- 11F0
         x"ff",  x"7f",  x"3f",  x"17",  x"13",  x"03",  x"03",  x"01", -- 11F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1200
         x"00",  x"04",  x"3f",  x"7b",  x"c1",  x"81",  x"00",  x"00", -- 1208
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"bf", -- 1210
         x"3f",  x"3f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1218
         x"ff",  x"e7",  x"ef",  x"f7",  x"ff",  x"ff",  x"ff",  x"ff", -- 1220
         x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f", -- 1228
         x"01",  x"29",  x"29",  x"29",  x"29",  x"29",  x"29",  x"29", -- 1230
         x"99",  x"c9",  x"e9",  x"c1",  x"99",  x"99",  x"99",  x"c1", -- 1238
         x"21",  x"2d",  x"2d",  x"2d",  x"0d",  x"2d",  x"2d",  x"21", -- 1240
         x"c3",  x"99",  x"99",  x"f9",  x"f1",  x"99",  x"99",  x"c3", -- 1248
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"9f",  x"9f", -- 1250
         x"99",  x"99",  x"99",  x"93",  x"8f",  x"95",  x"99",  x"99", -- 1258
         x"99",  x"89",  x"81",  x"91",  x"99",  x"99",  x"99",  x"99", -- 1260
         x"1e",  x"7c",  x"f8",  x"f0",  x"e0",  x"c1",  x"c7",  x"87", -- 1268
         x"c3",  x"99",  x"f9",  x"c1",  x"99",  x"99",  x"99",  x"c3", -- 1270
         x"c3",  x"99",  x"99",  x"99",  x"c3",  x"99",  x"99",  x"c3", -- 1278
         x"9f",  x"9f",  x"cf",  x"cf",  x"e7",  x"f3",  x"f9",  x"81", -- 1280
         x"c3",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"99",  x"c3", -- 1288
         x"81",  x"99",  x"f9",  x"f9",  x"83",  x"9f",  x"9f",  x"81", -- 1290
         x"f9",  x"f9",  x"f9",  x"c1",  x"99",  x"99",  x"99",  x"99", -- 1298
         x"c3",  x"99",  x"99",  x"f9",  x"f3",  x"99",  x"99",  x"c3", -- 12A0
         x"81",  x"9f",  x"cf",  x"e3",  x"f9",  x"99",  x"99",  x"c3", -- 12A8
         x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"c7",  x"e7", -- 12B0
         x"00",  x"99",  x"99",  x"99",  x"99",  x"99",  x"c9",  x"e1", -- 12B8
         x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"a5",  x"81", -- 12C0
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"99",  x"99", -- 12C8
         x"99",  x"99",  x"99",  x"81",  x"99",  x"99",  x"c9",  x"e1", -- 12D0
         x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"81", -- 12D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"81",  x"ff",  x"ff",  x"ff", -- 12E0
         x"c3",  x"99",  x"99",  x"f9",  x"81",  x"99",  x"99",  x"99", -- 12E8
         x"9f",  x"9f",  x"9f",  x"83",  x"99",  x"99",  x"99",  x"83", -- 12F0
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"99",  x"83", -- 12F8
         x"9f",  x"9f",  x"9f",  x"9f",  x"9f",  x"9f",  x"99",  x"83", -- 1300
         x"c3",  x"99",  x"99",  x"9f",  x"81",  x"99",  x"99",  x"c3", -- 1308
         x"99",  x"99",  x"99",  x"99",  x"81",  x"99",  x"99",  x"99", -- 1310
         x"c3",  x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"c3", -- 1318
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1320
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1328
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1330
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1338
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1340
         x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"c9",  x"e1", -- 1348
         x"29",  x"29",  x"29",  x"29",  x"01",  x"29",  x"29",  x"29", -- 1350
         x"83",  x"99",  x"99",  x"99",  x"83",  x"99",  x"99",  x"83", -- 1358
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"03",  x"ff", -- 1360
         x"e7",  x"ff",  x"f3",  x"ff",  x"ff",  x"ff",  x"fc",  x"ff", -- 1368
         x"0f",  x"ff",  x"f1",  x"ff",  x"ff",  x"ff",  x"f1",  x"ff", -- 1370
         x"80",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c4",  x"ff", -- 1378
         x"ff",  x"cf",  x"ff",  x"ff",  x"ff",  x"f3",  x"ff",  x"e0", -- 1380
         x"ff",  x"e3",  x"ff",  x"ff",  x"ff",  x"8f",  x"ff",  x"e7", -- 1388
         x"ff",  x"1f",  x"ff",  x"ff",  x"ff",  x"fb",  x"ff",  x"07", -- 1390
         x"ff",  x"c4",  x"ff",  x"ff",  x"ff",  x"c7",  x"ff",  x"80", -- 1398
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 13A0
         x"83",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c3",  x"ff", -- 13A8
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"1f",  x"1f", -- 13B0
         x"83",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c7",  x"ff", -- 13B8
         x"ff",  x"e7",  x"ff",  x"ff",  x"ff",  x"f1",  x"ff",  x"07", -- 13C0
         x"00",  x"28",  x"29",  x"29",  x"29",  x"29",  x"29",  x"29", -- 13C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fb",  x"ff",  x"07", -- 13D0
         x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c7",  x"ff",  x"80", -- 13D8
         x"1f",  x"ff",  x"f3",  x"ff",  x"ff",  x"ff",  x"f0",  x"ff", -- 13E0
         x"f8",  x"ff",  x"c3",  x"ff",  x"ff",  x"ff",  x"3c",  x"ff", -- 13E8
         x"c1",  x"ff",  x"e3",  x"ff",  x"ff",  x"ff",  x"e3",  x"ff", -- 13F0
         x"3c",  x"99",  x"99",  x"c3",  x"c3",  x"99",  x"99",  x"3c", -- 13F8
         x"ff",  x"07",  x"ff",  x"ff",  x"ff",  x"c3",  x"ff",  x"1f", -- 1400
         x"ff",  x"3c",  x"ff",  x"ff",  x"ff",  x"cf",  x"ff",  x"f8", -- 1408
         x"ff",  x"03",  x"ff",  x"ff",  x"ff",  x"e3",  x"ff",  x"c1", -- 1410
         x"ff",  x"c4",  x"ff",  x"ff",  x"ff",  x"07",  x"ff",  x"f3", -- 1418
         x"1f",  x"ff",  x"f3",  x"ff",  x"ff",  x"ff",  x"fc",  x"ff", -- 1420
         x"f8",  x"ff",  x"c3",  x"ff",  x"ff",  x"ff",  x"3f",  x"ff", -- 1428
         x"e0",  x"ff",  x"f1",  x"ff",  x"ff",  x"ff",  x"e7",  x"ff", -- 1430
         x"83",  x"ff",  x"c7",  x"ff",  x"ff",  x"ff",  x"c0",  x"ff", -- 1438
         x"ff",  x"fc",  x"ff",  x"ff",  x"ff",  x"c3",  x"ff",  x"1f", -- 1440
         x"ff",  x"3f",  x"ff",  x"ff",  x"ff",  x"cf",  x"ff",  x"f8", -- 1448
         x"ff",  x"9f",  x"ff",  x"ff",  x"ff",  x"f1",  x"ff",  x"e0", -- 1450
         x"ff",  x"c4",  x"ff",  x"ff",  x"ff",  x"07",  x"ff",  x"f3", -- 1458
         x"77",  x"1b",  x"0f",  x"01",  x"80",  x"f0",  x"e0",  x"c0", -- 1460
         x"e7",  x"81",  x"a5",  x"a5",  x"a5",  x"a5",  x"81",  x"e7", -- 1468
         x"cf",  x"cf",  x"ff",  x"cf",  x"cf",  x"cf",  x"cf",  x"cf", -- 1470
         x"01",  x"31",  x"33",  x"33",  x"33",  x"33",  x"33",  x"33", -- 1478
         x"ff",  x"ff",  x"fe",  x"fe",  x"fe",  x"f8",  x"00",  x"00", -- 1480
         x"c3",  x"99",  x"99",  x"9f",  x"9f",  x"99",  x"99",  x"c3", -- 1488
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00", -- 1490
         x"00",  x"03",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1498
         x"00",  x"00",  x"00",  x"1f",  x"1f",  x"7f",  x"ff",  x"ff", -- 14A0
         x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"1f",  x"00",  x"00", -- 14A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 14B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 14B8
         x"00",  x"00",  x"00",  x"f8",  x"fc",  x"ff",  x"ff",  x"ff", -- 14C0
         x"00",  x"80",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 14C8
         x"81",  x"e1",  x"f1",  x"f3",  x"3f",  x"ff",  x"7f",  x"ff", -- 14D0
         x"03",  x"0f",  x"1f",  x"9e",  x"f8",  x"ff",  x"fd",  x"ff", -- 14D8
         x"ff",  x"b7",  x"f7",  x"f3",  x"a3",  x"07",  x"0f",  x"1f", -- 14E0
         x"ff",  x"dd",  x"df",  x"9f",  x"8b",  x"ce",  x"e4",  x"f8", -- 14E8
         x"01",  x"00",  x"40",  x"04",  x"00",  x"10",  x"02",  x"00", -- 14F0
         x"80",  x"c0",  x"c0",  x"e0",  x"4c",  x"0c",  x"06",  x"ff", -- 14F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1500
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1508
         x"f8",  x"e0",  x"e0",  x"e3",  x"83",  x"87",  x"1e",  x"1c", -- 1510
         x"ff",  x"ff",  x"f1",  x"80",  x"80",  x"08",  x"1c",  x"3e", -- 1518
         x"fe",  x"f8",  x"e0",  x"80",  x"00",  x"00",  x"00",  x"00", -- 1520
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"f8",  x"e0",  x"80", -- 1528
         x"03",  x"03",  x"71",  x"f1",  x"f0",  x"70",  x"00",  x"ff", -- 1530
         x"80",  x"80",  x"80",  x"90",  x"10",  x"38",  x"fe",  x"98", -- 1538
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1540
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1548
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1550
         x"2f",  x"6f",  x"7f",  x"df",  x"df",  x"4f",  x"6f",  x"0f", -- 1558
         x"78",  x"34",  x"14",  x"18",  x"34",  x"64",  x"64",  x"74", -- 1560
         x"5f",  x"5f",  x"3f",  x"3f",  x"5f",  x"0f",  x"af",  x"af", -- 1568
         x"78",  x"60",  x"2c",  x"3e",  x"1a",  x"32",  x"52",  x"50", -- 1570
         x"39",  x"29",  x"29",  x"01",  x"01",  x"11",  x"39",  x"7d", -- 1578
         x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"1f",  x"07",  x"01", -- 1580
         x"7f",  x"1f",  x"07",  x"01",  x"00",  x"00",  x"00",  x"00", -- 1588
         x"ff",  x"e7",  x"c1",  x"80",  x"00",  x"00",  x"18",  x"3c", -- 1590
         x"ff",  x"7f",  x"3f",  x"1f",  x"0f",  x"07",  x"03",  x"01", -- 1598
         x"ff",  x"7f",  x"1f",  x"07",  x"01",  x"00",  x"00",  x"00", -- 15A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7c",  x"38",  x"00", -- 15A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15B0
         x"3c",  x"0f",  x"07",  x"03",  x"00",  x"00",  x"00",  x"00", -- 15B8
         x"f0",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00",  x"00", -- 15C0
         x"90",  x"f8",  x"c0",  x"80",  x"99",  x"0f",  x"1f",  x"3f", -- 15C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"e0",  x"f8", -- 15D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15D8
         x"03",  x"07",  x"07",  x"0f",  x"0c",  x"00",  x"00",  x"00", -- 15E0
         x"00",  x"00",  x"00",  x"1c",  x"3e",  x"3f",  x"ed",  x"f3", -- 15E8
         x"00",  x"00",  x"00",  x"00",  x"04",  x"0e",  x"0f",  x"1f", -- 15F0
         x"00",  x"00",  x"00",  x"1c",  x"bc",  x"f9",  x"f3",  x"ff", -- 15F8
         x"ff",  x"fc",  x"f0",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 1600
         x"ff",  x"fe",  x"fc",  x"f8",  x"f0",  x"e0",  x"c0",  x"80", -- 1608
         x"ff",  x"ff",  x"e3",  x"80",  x"00",  x"00",  x"00",  x"00", -- 1610
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1618
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1620
         x"e3",  x"c1",  x"80",  x"08",  x"1c",  x"ff",  x"fb",  x"fc", -- 1628
         x"f0",  x"e0",  x"e0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 1630
         x"00",  x"00",  x"00",  x"08",  x"1c",  x"78",  x"f0",  x"e0", -- 1638
         x"f9",  x"f0",  x"c0",  x"c0",  x"81",  x"03",  x"1f",  x"0e", -- 1640
         x"80",  x"c0",  x"f0",  x"f0",  x"f8",  x"fc",  x"7f",  x"3f", -- 1648
         x"ff",  x"ff",  x"ff",  x"ff",  x"9f",  x"83",  x"80",  x"00", -- 1650
         x"80",  x"e0",  x"e0",  x"f0",  x"f8",  x"f8",  x"fc",  x"fe", -- 1658
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1660
         x"ff",  x"ff",  x"33",  x"01",  x"00",  x"90",  x"f0",  x"f8", -- 1668
         x"af",  x"df",  x"fe",  x"78",  x"19",  x"03",  x"03",  x"1f", -- 1670
         x"ff",  x"f8",  x"e0",  x"c0",  x"80",  x"83",  x"07",  x"03", -- 1678
         x"ff",  x"dd",  x"0c",  x"07",  x"01",  x"00",  x"00",  x"00", -- 1680
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1688
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1690
         x"c0",  x"82",  x"0e",  x"0e",  x"1e",  x"8f",  x"87",  x"c1", -- 1698
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"e3",  x"c0",  x"81", -- 16A0
         x"7f",  x"1f",  x"07",  x"3f",  x"0f",  x"03",  x"01",  x"00", -- 16A8
         x"c3",  x"81",  x"80",  x"0c",  x"1e",  x"b7",  x"e9",  x"fd", -- 16B0
         x"81",  x"e0",  x"f0",  x"f0",  x"fc",  x"fe",  x"fe",  x"ff", -- 16B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 16C0
         x"00",  x"00",  x"00",  x"80",  x"80",  x"80",  x"00",  x"00", -- 16C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16D8
         x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe", -- 16E0
         x"07",  x"83",  x"41",  x"c3",  x"e3",  x"e3",  x"f1",  x"fc", -- 16E8
         x"7f",  x"7f",  x"fb",  x"fd",  x"f0",  x"f9",  x"e3",  x"ff", -- 16F0
         x"ff",  x"ff",  x"cf",  x"c7",  x"83",  x"83",  x"c1",  x"e1", -- 16F8
         x"ff",  x"ff",  x"f6",  x"e0",  x"fc",  x"f8",  x"f0",  x"f0", -- 1700
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1708
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1710
         x"e0",  x"40",  x"40",  x"40",  x"40",  x"00",  x"00",  x"00", -- 1718
         x"ff",  x"77",  x"32",  x"22",  x"22",  x"02",  x"00",  x"00", -- 1720
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1728
         x"1f",  x"07",  x"03",  x"03",  x"e3",  x"61",  x"70",  x"f8", -- 1730
         x"05",  x"43",  x"63",  x"f1",  x"f1",  x"c1",  x"03",  x"07", -- 1738
         x"d0",  x"5c",  x"b8",  x"f9",  x"e1",  x"83",  x"0f",  x"1e", -- 1740
         x"7c",  x"ec",  x"c0",  x"81",  x"93",  x"0f",  x"0e",  x"3c", -- 1748
         x"3c",  x"31",  x"7d",  x"ee",  x"d3",  x"f9",  x"69",  x"1c", -- 1750
         x"13",  x"01",  x"81",  x"80",  x"c8",  x"78",  x"58",  x"3e", -- 1758
         x"e1",  x"c1",  x"83",  x"c3",  x"c7",  x"01",  x"60",  x"b8", -- 1760
         x"df",  x"3e",  x"f4",  x"c0",  x"80",  x"13",  x"1f",  x"3f", -- 1768
         x"79",  x"1e",  x"0f",  x"01",  x"80",  x"f0",  x"f8",  x"fc", -- 1770
         x"73",  x"79",  x"ec",  x"c0",  x"80",  x"01",  x"13",  x"3f", -- 1778
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1780
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1788
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1790
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1798
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1800
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1808
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1810
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1818
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1820
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1828
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80", -- 1830
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80", -- 1838
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 1840
         x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"80",  x"ff", -- 1848
         x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1850
         x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1858
         x"80",  x"80",  x"80",  x"88",  x"80",  x"80",  x"80",  x"ff", -- 1860
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1868
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1870
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1878
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1880
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1888
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1890
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1898
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18D0
         x"01",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe", -- 18D8
         x"c0",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf", -- 18E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 18E8
         x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"01", -- 18F0
         x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"bf",  x"c0", -- 18F8
         x"fa",  x"f7",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1900
         x"bf",  x"df",  x"ef",  x"7f",  x"7f",  x"ff",  x"ff",  x"ff", -- 1908
         x"ff",  x"f0",  x"f9",  x"fd",  x"fd",  x"ff",  x"ff",  x"ff", -- 1910
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"7f",  x"5f",  x"bf", -- 1918
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"f8",  x"f0",  x"c0", -- 1920
         x"ff",  x"ff",  x"7f",  x"7f",  x"3f",  x"1f",  x"0f",  x"03", -- 1928
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"f8",  x"f0",  x"c0", -- 1930
         x"ff",  x"ff",  x"7f",  x"7f",  x"3f",  x"1f",  x"0f",  x"03", -- 1938
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1940
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1948
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1950
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1958
         x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"f8",  x"f0",  x"c0", -- 1960
         x"ff",  x"ff",  x"7f",  x"7f",  x"3f",  x"1f",  x"0f",  x"03", -- 1968
         x"7f",  x"7f",  x"7f",  x"0f",  x"e7",  x"e7",  x"e7",  x"00", -- 1970
         x"7e",  x"7e",  x"7e",  x"00",  x"e7",  x"e7",  x"e7",  x"00", -- 1978
         x"00",  x"00",  x"00",  x"1c",  x"00",  x"00",  x"00",  x"00", -- 1980
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1988
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1990
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1998
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19A8
         x"fe",  x"fe",  x"fe",  x"f0",  x"f7",  x"f7",  x"f7",  x"00", -- 19B0
         x"00",  x"00",  x"00",  x"00",  x"18",  x"18",  x"3c",  x"7e", -- 19B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19C0
         x"7e",  x"02",  x"02",  x"00",  x"e7",  x"20",  x"20",  x"00", -- 19C8
         x"88",  x"c0",  x"80",  x"80",  x"80",  x"00",  x"00",  x"00", -- 19D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19E8
         x"00",  x"00",  x"02",  x"07",  x"27",  x"7f",  x"7f",  x"7f", -- 19F0
         x"00",  x"80",  x"c0",  x"e8",  x"ec",  x"fc",  x"fc",  x"fe", -- 19F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A00
         x"ff",  x"fb",  x"c0",  x"84",  x"3e",  x"7e",  x"ff",  x"ff", -- 1A08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"bf", -- 1A10
         x"3f",  x"3f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A18
         x"ff",  x"e7",  x"ef",  x"f7",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A20
         x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f", -- 1A28
         x"01",  x"29",  x"29",  x"29",  x"29",  x"29",  x"29",  x"29", -- 1A30
         x"99",  x"c9",  x"e9",  x"c1",  x"99",  x"99",  x"99",  x"c1", -- 1A38
         x"21",  x"2d",  x"2d",  x"2d",  x"0d",  x"2d",  x"2d",  x"21", -- 1A40
         x"c3",  x"99",  x"99",  x"f9",  x"f1",  x"99",  x"99",  x"c3", -- 1A48
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"9f",  x"9f", -- 1A50
         x"99",  x"99",  x"99",  x"93",  x"8f",  x"95",  x"99",  x"99", -- 1A58
         x"99",  x"89",  x"81",  x"91",  x"99",  x"99",  x"99",  x"99", -- 1A60
         x"e1",  x"83",  x"07",  x"0f",  x"1f",  x"3e",  x"38",  x"78", -- 1A68
         x"c3",  x"99",  x"f9",  x"c1",  x"99",  x"99",  x"99",  x"c3", -- 1A70
         x"c3",  x"99",  x"99",  x"99",  x"c3",  x"99",  x"99",  x"c3", -- 1A78
         x"9f",  x"9f",  x"cf",  x"cf",  x"e7",  x"f3",  x"f9",  x"81", -- 1A80
         x"c3",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"99",  x"c3", -- 1A88
         x"81",  x"99",  x"f9",  x"f9",  x"83",  x"9f",  x"9f",  x"81", -- 1A90
         x"f9",  x"f9",  x"f9",  x"c1",  x"99",  x"99",  x"99",  x"99", -- 1A98
         x"c3",  x"99",  x"99",  x"f9",  x"f3",  x"99",  x"99",  x"c3", -- 1AA0
         x"81",  x"9f",  x"cf",  x"e3",  x"f9",  x"99",  x"99",  x"c3", -- 1AA8
         x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"c7",  x"e7", -- 1AB0
         x"00",  x"99",  x"99",  x"99",  x"99",  x"99",  x"c9",  x"e1", -- 1AB8
         x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"a5",  x"81", -- 1AC0
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"99",  x"99", -- 1AC8
         x"99",  x"99",  x"99",  x"81",  x"99",  x"99",  x"c9",  x"e1", -- 1AD0
         x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"81", -- 1AD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"81",  x"ff",  x"ff",  x"ff", -- 1AE0
         x"c3",  x"99",  x"99",  x"f9",  x"81",  x"99",  x"99",  x"99", -- 1AE8
         x"9f",  x"9f",  x"9f",  x"83",  x"99",  x"99",  x"99",  x"83", -- 1AF0
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"99",  x"83", -- 1AF8
         x"9f",  x"9f",  x"9f",  x"9f",  x"9f",  x"9f",  x"99",  x"83", -- 1B00
         x"c3",  x"99",  x"99",  x"9f",  x"81",  x"99",  x"99",  x"c3", -- 1B08
         x"99",  x"99",  x"99",  x"99",  x"81",  x"99",  x"99",  x"99", -- 1B10
         x"c3",  x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"c3", -- 1B18
         x"00",  x"00",  x"80",  x"a0",  x"e0",  x"e8",  x"f8",  x"fe", -- 1B20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B40
         x"99",  x"99",  x"99",  x"99",  x"99",  x"99",  x"c9",  x"e1", -- 1B48
         x"29",  x"29",  x"29",  x"29",  x"01",  x"29",  x"29",  x"29", -- 1B50
         x"83",  x"99",  x"99",  x"99",  x"83",  x"99",  x"99",  x"83", -- 1B58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B60
         x"ff",  x"f7",  x"f3",  x"f9",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B68
         x"ff",  x"e3",  x"f1",  x"f1",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B70
         x"ff",  x"c3",  x"c7",  x"c7",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B78
         x"ff",  x"ff",  x"ff",  x"ff",  x"f3",  x"f3",  x"f1",  x"ff", -- 1B80
         x"ff",  x"ff",  x"ff",  x"ff",  x"07",  x"8f",  x"cf",  x"ff", -- 1B88
         x"ff",  x"ff",  x"ff",  x"ff",  x"fd",  x"fb",  x"e3",  x"ff", -- 1B90
         x"ff",  x"ff",  x"ff",  x"ff",  x"c7",  x"c7",  x"c3",  x"ff", -- 1B98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1BA0
         x"ff",  x"c7",  x"c7",  x"c7",  x"ff",  x"ff",  x"ff",  x"ff", -- 1BA8
         x"83",  x"99",  x"99",  x"99",  x"83",  x"9f",  x"1f",  x"1f", -- 1BB0
         x"ff",  x"c7",  x"c7",  x"c7",  x"ff",  x"ff",  x"ff",  x"ff", -- 1BB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"f1",  x"f1",  x"e1",  x"ff", -- 1BC0
         x"00",  x"28",  x"29",  x"29",  x"29",  x"29",  x"29",  x"29", -- 1BC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"fd",  x"fb",  x"e3",  x"ff", -- 1BD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"c7",  x"c7",  x"c3",  x"ff", -- 1BD8
         x"ff",  x"07",  x"f3",  x"f9",  x"ff",  x"ff",  x"ff",  x"ff", -- 1BE0
         x"ff",  x"e0",  x"c3",  x"87",  x"ff",  x"ff",  x"ff",  x"ff", -- 1BE8
         x"ff",  x"e3",  x"e3",  x"e3",  x"ff",  x"ff",  x"ff",  x"ff", -- 1BF0
         x"3c",  x"99",  x"99",  x"c3",  x"c3",  x"99",  x"99",  x"3c", -- 1BF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"e1",  x"c3",  x"0f",  x"ff", -- 1C00
         x"ff",  x"ff",  x"ff",  x"ff",  x"9f",  x"cf",  x"e0",  x"ff", -- 1C08
         x"ff",  x"ff",  x"ff",  x"ff",  x"e3",  x"e3",  x"e3",  x"ff", -- 1C10
         x"ff",  x"ff",  x"ff",  x"ff",  x"c7",  x"07",  x"c7",  x"ff", -- 1C18
         x"ff",  x"07",  x"f3",  x"f9",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C20
         x"ff",  x"e0",  x"c3",  x"87",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C28
         x"ff",  x"f1",  x"f1",  x"e3",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C30
         x"ff",  x"c7",  x"c7",  x"c7",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C38
         x"ff",  x"ff",  x"ff",  x"ff",  x"e1",  x"c3",  x"07",  x"ff", -- 1C40
         x"ff",  x"ff",  x"ff",  x"ff",  x"9f",  x"cf",  x"e0",  x"ff", -- 1C48
         x"ff",  x"ff",  x"ff",  x"ff",  x"f1",  x"f1",  x"f0",  x"ff", -- 1C50
         x"ff",  x"ff",  x"ff",  x"ff",  x"c7",  x"07",  x"c7",  x"ff", -- 1C58
         x"88",  x"e4",  x"f0",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C60
         x"e7",  x"81",  x"a5",  x"a5",  x"a5",  x"a5",  x"81",  x"e7", -- 1C68
         x"cf",  x"cf",  x"ff",  x"cf",  x"cf",  x"cf",  x"cf",  x"cf", -- 1C70
         x"01",  x"31",  x"33",  x"33",  x"33",  x"33",  x"33",  x"33", -- 1C78
         x"ff",  x"ff",  x"fe",  x"fe",  x"fe",  x"f8",  x"00",  x"00", -- 1C80
         x"c3",  x"99",  x"99",  x"9f",  x"9f",  x"99",  x"99",  x"c3", -- 1C88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00", -- 1C90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1CA0
         x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"1f",  x"00",  x"00", -- 1CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1CB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1CC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1CC8
         x"81",  x"e1",  x"f1",  x"f3",  x"3f",  x"ff",  x"ff",  x"ff", -- 1CD0
         x"03",  x"0f",  x"1f",  x"9e",  x"f8",  x"ff",  x"ff",  x"ff", -- 1CD8
         x"ff",  x"f7",  x"f7",  x"f3",  x"a3",  x"07",  x"0f",  x"1f", -- 1CE0
         x"ff",  x"df",  x"df",  x"9f",  x"8b",  x"ce",  x"e4",  x"f8", -- 1CE8
         x"fe",  x"ff",  x"bf",  x"fb",  x"ff",  x"ef",  x"fd",  x"ff", -- 1CF0
         x"1f",  x"0f",  x"0f",  x"1f",  x"b1",  x"f0",  x"f9",  x"00", -- 1CF8
         x"00",  x"80",  x"c1",  x"c1",  x"c3",  x"e3",  x"e3",  x"f7", -- 1D00
         x"01",  x"07",  x"01",  x"03",  x"07",  x"03",  x"07",  x"0f", -- 1D08
         x"07",  x"1f",  x"1f",  x"1c",  x"7c",  x"78",  x"e1",  x"e3", -- 1D10
         x"00",  x"00",  x"0e",  x"7f",  x"7f",  x"f7",  x"e3",  x"c1", -- 1D18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D28
         x"fc",  x"fc",  x"86",  x"02",  x"03",  x"87",  x"ff",  x"00", -- 1D30
         x"7f",  x"7f",  x"7f",  x"6f",  x"ef",  x"c7",  x"01",  x"67", -- 1D38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D48
         x"ff",  x"75",  x"a5",  x"14",  x"02",  x"00",  x"00",  x"b9", -- 1D50
         x"d0",  x"90",  x"80",  x"20",  x"20",  x"b0",  x"90",  x"f0", -- 1D58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D60
         x"a0",  x"a0",  x"c0",  x"c0",  x"a0",  x"f0",  x"50",  x"50", -- 1D68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D70
         x"39",  x"29",  x"29",  x"01",  x"01",  x"11",  x"39",  x"7d", -- 1D78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D88
         x"00",  x"18",  x"3e",  x"7f",  x"ff",  x"ff",  x"e7",  x"c3", -- 1D90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DA8
         x"07",  x"8f",  x"9f",  x"df",  x"df",  x"df",  x"df",  x"ff", -- 1DB0
         x"c3",  x"f0",  x"f8",  x"fc",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DB8
         x"0f",  x"3f",  x"3f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DC0
         x"6f",  x"07",  x"3f",  x"7f",  x"66",  x"f0",  x"e0",  x"c0", -- 1DC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"1f",  x"07", -- 1DD0
         x"00",  x"8c",  x"d8",  x"dc",  x"fe",  x"fc",  x"fe",  x"ff", -- 1DD8
         x"fc",  x"f8",  x"f8",  x"f0",  x"f3",  x"ff",  x"ff",  x"ff", -- 1DE0
         x"ff",  x"ff",  x"ff",  x"e3",  x"c1",  x"c0",  x"12",  x"0c", -- 1DE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"fb",  x"f1",  x"f0",  x"e0", -- 1DF0
         x"ff",  x"ff",  x"ff",  x"e3",  x"43",  x"06",  x"0c",  x"00", -- 1DF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E08
         x"00",  x"00",  x"1c",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E20
         x"1c",  x"3e",  x"7f",  x"f7",  x"e3",  x"00",  x"04",  x"03", -- 1E28
         x"0f",  x"1f",  x"1f",  x"3f",  x"7f",  x"ff",  x"ff",  x"ff", -- 1E30
         x"ff",  x"ff",  x"ff",  x"f7",  x"e3",  x"87",  x"0f",  x"1f", -- 1E38
         x"06",  x"0f",  x"3f",  x"3f",  x"7e",  x"fc",  x"e0",  x"f1", -- 1E40
         x"7f",  x"3f",  x"0f",  x"0f",  x"07",  x"03",  x"80",  x"c0", -- 1E48
         x"00",  x"00",  x"00",  x"00",  x"60",  x"7c",  x"7f",  x"ff", -- 1E50
         x"7f",  x"1f",  x"1f",  x"0f",  x"07",  x"07",  x"03",  x"01", -- 1E58
         x"00",  x"00",  x"80",  x"e0",  x"00",  x"c0",  x"f0",  x"c0", -- 1E60
         x"00",  x"00",  x"cc",  x"fe",  x"ff",  x"6f",  x"0f",  x"07", -- 1E68
         x"50",  x"20",  x"01",  x"87",  x"e6",  x"fc",  x"fc",  x"e0", -- 1E70
         x"00",  x"07",  x"1f",  x"3f",  x"7f",  x"7c",  x"f8",  x"fc", -- 1E78
         x"00",  x"22",  x"f3",  x"f8",  x"fe",  x"ff",  x"ff",  x"ff", -- 1E80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E90
         x"3f",  x"7d",  x"f1",  x"f1",  x"e1",  x"70",  x"78",  x"3e", -- 1E98
         x"e0",  x"f0",  x"c0",  x"fc",  x"f0",  x"fc",  x"ff",  x"fe", -- 1EA0
         x"80",  x"e0",  x"f8",  x"c0",  x"f0",  x"fc",  x"fe",  x"ff", -- 1EA8
         x"3c",  x"7e",  x"7f",  x"f3",  x"e1",  x"48",  x"16",  x"02", -- 1EB0
         x"7e",  x"1f",  x"0f",  x"0f",  x"03",  x"01",  x"01",  x"00", -- 1EB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1EC0
         x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f",  x"ff",  x"ff", -- 1EC8
         x"00",  x"80",  x"e0",  x"c0",  x"f8",  x"e0",  x"fc",  x"fe", -- 1ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"04",  x"0e", -- 1ED8
         x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01", -- 1EE0
         x"f8",  x"7c",  x"be",  x"3c",  x"1c",  x"1c",  x"8e",  x"e3", -- 1EE8
         x"80",  x"80",  x"04",  x"02",  x"0f",  x"06",  x"1c",  x"00", -- 1EF0
         x"f0",  x"38",  x"3c",  x"3e",  x"7f",  x"7f",  x"3f",  x"1f", -- 1EF8
         x"00",  x"00",  x"09",  x"1f",  x"03",  x"07",  x"0f",  x"0f", -- 1F00
         x"00",  x"10",  x"b8",  x"fe",  x"f0",  x"fc",  x"fe",  x"fe", -- 1F08
         x"1f",  x"3f",  x"1f",  x"3f",  x"7f",  x"7f",  x"ff",  x"ff", -- 1F10
         x"1f",  x"bf",  x"bf",  x"bf",  x"bf",  x"ff",  x"ff",  x"ff", -- 1F18
         x"00",  x"88",  x"cd",  x"dd",  x"dd",  x"fd",  x"ff",  x"ff", -- 1F20
         x"03",  x"01",  x"01",  x"03",  x"07",  x"3f",  x"1f",  x"3f", -- 1F28
         x"e0",  x"f8",  x"fc",  x"fc",  x"1c",  x"9e",  x"8f",  x"07", -- 1F30
         x"fa",  x"bc",  x"9c",  x"0e",  x"0e",  x"3e",  x"fc",  x"f8", -- 1F38
         x"2f",  x"a3",  x"47",  x"06",  x"1e",  x"7c",  x"f0",  x"e1", -- 1F40
         x"83",  x"13",  x"3f",  x"7e",  x"6c",  x"f0",  x"f1",  x"c3", -- 1F48
         x"c3",  x"ce",  x"82",  x"11",  x"2c",  x"06",  x"96",  x"e3", -- 1F50
         x"ec",  x"fe",  x"7e",  x"7f",  x"37",  x"87",  x"a7",  x"c1", -- 1F58
         x"1e",  x"3e",  x"7c",  x"3c",  x"38",  x"fe",  x"9f",  x"47", -- 1F60
         x"20",  x"c1",  x"0b",  x"3f",  x"7f",  x"ec",  x"e0",  x"c0", -- 1F68
         x"86",  x"e1",  x"f0",  x"fe",  x"7f",  x"0f",  x"07",  x"03", -- 1F70
         x"8c",  x"86",  x"13",  x"3f",  x"7f",  x"fe",  x"ec",  x"c0", -- 1F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
