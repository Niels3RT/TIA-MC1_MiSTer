library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_g2 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_g2;

architecture rtl of rom_g2 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"f0",  x"21",  x"ad",  x"16",  x"11",  x"89",  x"f1",  x"cd", -- 0000
         x"4d",  x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"ff",  x"f0", -- 0008
         x"af",  x"32",  x"00",  x"f1",  x"32",  x"87",  x"f1",  x"22", -- 0010
         x"03",  x"f1",  x"c3",  x"91",  x"1f",  x"af",  x"32",  x"0a", -- 0018
         x"f1",  x"32",  x"eb",  x"f0",  x"21",  x"87",  x"f1",  x"22", -- 0020
         x"14",  x"f0",  x"21",  x"77",  x"f1",  x"22",  x"17",  x"f0", -- 0028
         x"21",  x"b5",  x"16",  x"11",  x"87",  x"f1",  x"cd",  x"4d", -- 0030
         x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"00",  x"f1",  x"3e", -- 0038
         x"07",  x"32",  x"f7",  x"f0",  x"32",  x"f5",  x"f0",  x"32", -- 0040
         x"f8",  x"f0",  x"21",  x"ee",  x"16",  x"22",  x"03",  x"f1", -- 0048
         x"3e",  x"01",  x"32",  x"ed",  x"f0",  x"c9",  x"af",  x"32", -- 0050
         x"8a",  x"f1",  x"32",  x"a6",  x"f1",  x"32",  x"14",  x"f1", -- 0058
         x"32",  x"1a",  x"f1",  x"32",  x"f5",  x"f0",  x"32",  x"f8", -- 0060
         x"f0",  x"32",  x"e9",  x"f0",  x"32",  x"eb",  x"f0",  x"cd", -- 0068
         x"e3",  x"0f",  x"3e",  x"01",  x"32",  x"19",  x"f1",  x"32", -- 0070
         x"e8",  x"f0",  x"3e",  x"bf",  x"32",  x"27",  x"f0",  x"32", -- 0078
         x"21",  x"f0",  x"3e",  x"a7",  x"32",  x"24",  x"f0",  x"3e", -- 0080
         x"a7",  x"32",  x"5f",  x"f1",  x"32",  x"60",  x"f1",  x"c6", -- 0088
         x"10",  x"32",  x"61",  x"f1",  x"32",  x"62",  x"f1",  x"af", -- 0090
         x"32",  x"6f",  x"f1",  x"32",  x"71",  x"f1",  x"c6",  x"10", -- 0098
         x"32",  x"70",  x"f1",  x"32",  x"72",  x"f1",  x"21",  x"29", -- 00A0
         x"f0",  x"11",  x"7f",  x"f1",  x"cd",  x"4d",  x"1b",  x"3a", -- 00A8
         x"f9",  x"f0",  x"32",  x"fa",  x"f0",  x"c9",  x"db",  x"d2", -- 00B0
         x"e6",  x"20",  x"ca",  x"c2",  x"20",  x"3e",  x"59",  x"c3", -- 00B8
         x"fe",  x"20",  x"db",  x"d0",  x"47",  x"e6",  x"02",  x"ca", -- 00C0
         x"cf",  x"20",  x"3e",  x"47",  x"c3",  x"fe",  x"20",  x"78", -- 00C8
         x"e6",  x"20",  x"ca",  x"da",  x"20",  x"3e",  x"42",  x"c3", -- 00D0
         x"fe",  x"20",  x"db",  x"d1",  x"47",  x"e6",  x"02",  x"ca", -- 00D8
         x"e7",  x"20",  x"3e",  x"4a",  x"c3",  x"fe",  x"20",  x"78", -- 00E0
         x"e6",  x"20",  x"ca",  x"f2",  x"20",  x"3e",  x"4c",  x"c3", -- 00E8
         x"fe",  x"20",  x"3e",  x"53",  x"47",  x"3a",  x"a6",  x"f1", -- 00F0
         x"fe",  x"52",  x"ca",  x"fe",  x"20",  x"78",  x"47",  x"3a", -- 00F8
         x"a6",  x"f1",  x"b8",  x"78",  x"c2",  x"09",  x"21",  x"af", -- 0100
         x"c9",  x"b7",  x"f5",  x"cd",  x"e3",  x"0f",  x"f1",  x"c9", -- 0108
         x"3e",  x"68",  x"32",  x"84",  x"f1",  x"3e",  x"a5",  x"32", -- 0110
         x"64",  x"f1",  x"3e",  x"05",  x"32",  x"94",  x"f1",  x"c9", -- 0118
         x"01",  x"8b",  x"f1",  x"21",  x"9a",  x"f1",  x"3e",  x"05", -- 0120
         x"cd",  x"6d",  x"12",  x"01",  x"5b",  x"f1",  x"21",  x"8a", -- 0128
         x"f1",  x"af",  x"cd",  x"6d",  x"12",  x"c9",  x"cd",  x"20", -- 0130
         x"21",  x"32",  x"a4",  x"f1",  x"32",  x"a6",  x"f1",  x"32", -- 0138
         x"9c",  x"f1",  x"32",  x"15",  x"f1",  x"32",  x"16",  x"f1", -- 0140
         x"3e",  x"46",  x"32",  x"fa",  x"f0",  x"3e",  x"01",  x"32", -- 0148
         x"9b",  x"f1",  x"32",  x"13",  x"f1",  x"32",  x"14",  x"f1", -- 0150
         x"32",  x"19",  x"f1",  x"32",  x"a5",  x"f1",  x"32",  x"f6", -- 0158
         x"f0",  x"32",  x"f5",  x"f0",  x"32",  x"0e",  x"f1",  x"32", -- 0160
         x"0f",  x"f1",  x"32",  x"fb",  x"f0",  x"3c",  x"32",  x"fd", -- 0168
         x"f0",  x"3c",  x"32",  x"fc",  x"f0",  x"c9",  x"3e",  x"04", -- 0170
         x"11",  x"9a",  x"f1",  x"12",  x"1b",  x"05",  x"c2",  x"7b", -- 0178
         x"21",  x"cd",  x"9f",  x"1a",  x"c9",  x"21",  x"6b",  x"f1", -- 0180
         x"36",  x"03",  x"23",  x"36",  x"13",  x"23",  x"36",  x"03", -- 0188
         x"23",  x"36",  x"13",  x"23",  x"c9",  x"01",  x"5b",  x"f1", -- 0190
         x"3e",  x"95",  x"02",  x"03",  x"02",  x"03",  x"3e",  x"a5", -- 0198
         x"02",  x"03",  x"02",  x"03",  x"c9",  x"21",  x"7b",  x"f1", -- 01A0
         x"36",  x"d8",  x"23",  x"36",  x"00",  x"23",  x"36",  x"e8", -- 01A8
         x"23",  x"36",  x"f8",  x"23",  x"c9",  x"cd",  x"20",  x"21", -- 01B0
         x"cd",  x"95",  x"21",  x"21",  x"70",  x"17",  x"cd",  x"f8", -- 01B8
         x"21",  x"c3",  x"4c",  x"39",  x"cd",  x"20",  x"21",  x"21", -- 01C0
         x"30",  x"30",  x"22",  x"5b",  x"f1",  x"21",  x"40",  x"40", -- 01C8
         x"22",  x"5d",  x"f1",  x"c3",  x"dc",  x"21",  x"cd",  x"20", -- 01D0
         x"21",  x"cd",  x"95",  x"21",  x"21",  x"6c",  x"16",  x"cd", -- 01D8
         x"f8",  x"21",  x"c3",  x"4c",  x"39",  x"3a",  x"6b",  x"f1", -- 01E0
         x"fe",  x"c8",  x"d2",  x"f3",  x"21",  x"cd",  x"9f",  x"1a", -- 01E8
         x"c3",  x"4c",  x"39",  x"af",  x"32",  x"a4",  x"f1",  x"c9", -- 01F0
         x"11",  x"7b",  x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"15", -- 01F8
         x"f1",  x"cd",  x"85",  x"21",  x"3e",  x"01",  x"32",  x"a4", -- 0200
         x"f1",  x"3e",  x"0a",  x"32",  x"f5",  x"f0",  x"af",  x"32", -- 0208
         x"13",  x"f1",  x"c9",  x"21",  x"7f",  x"f1",  x"22",  x"08", -- 0210
         x"f0",  x"01",  x"30",  x"06",  x"cd",  x"20",  x"22",  x"c9", -- 0218
         x"21",  x"9e",  x"f1",  x"79",  x"86",  x"77",  x"23",  x"05", -- 0220
         x"c2",  x"23",  x"22",  x"c9",  x"21",  x"9e",  x"f1",  x"36", -- 0228
         x"35",  x"23",  x"36",  x"38",  x"23",  x"36",  x"3c",  x"23", -- 0230
         x"36",  x"4a",  x"23",  x"36",  x"50",  x"23",  x"36",  x"58", -- 0238
         x"c9",  x"0e",  x"30",  x"79",  x"cd",  x"9f",  x"1a",  x"0d", -- 0240
         x"c2",  x"44",  x"22",  x"c9",  x"3e",  x"4e",  x"77",  x"23", -- 0248
         x"3e",  x"76",  x"77",  x"3e",  x"e0",  x"32",  x"72",  x"f1", -- 0250
         x"c6",  x"08",  x"32",  x"73",  x"f1",  x"3e",  x"20",  x"32", -- 0258
         x"62",  x"f1",  x"c6",  x"06",  x"32",  x"63",  x"f1",  x"3e", -- 0260
         x"09",  x"32",  x"92",  x"f1",  x"21",  x"23",  x"17",  x"22", -- 0268
         x"a7",  x"f1",  x"21",  x"e0",  x"17",  x"22",  x"06",  x"f1", -- 0270
         x"3a",  x"a3",  x"f0",  x"86",  x"32",  x"e7",  x"f0",  x"c9", -- 0278
         x"cd",  x"36",  x"21",  x"21",  x"81",  x"f1",  x"22",  x"08", -- 0280
         x"f0",  x"3e",  x"03",  x"32",  x"1a",  x"f1",  x"cd",  x"85", -- 0288
         x"21",  x"36",  x"c0",  x"23",  x"36",  x"90",  x"23",  x"36", -- 0290
         x"40",  x"cd",  x"95",  x"21",  x"3e",  x"a5",  x"02",  x"03", -- 0298
         x"02",  x"03",  x"02",  x"cd",  x"a5",  x"21",  x"3a",  x"ff", -- 02A0
         x"f0",  x"77",  x"23",  x"77",  x"23",  x"77",  x"c9",  x"21", -- 02A8
         x"9e",  x"f1",  x"36",  x"3c",  x"23",  x"36",  x"40",  x"23", -- 02B0
         x"36",  x"45",  x"23",  x"36",  x"42",  x"23",  x"36",  x"48", -- 02B8
         x"23",  x"36",  x"50",  x"c9",  x"3a",  x"6b",  x"f1",  x"c6", -- 02C0
         x"08",  x"32",  x"6b",  x"f1",  x"3a",  x"5b",  x"f1",  x"c6", -- 02C8
         x"08",  x"32",  x"5b",  x"f1",  x"af",  x"32",  x"13",  x"f1", -- 02D0
         x"32",  x"14",  x"f1",  x"32",  x"8a",  x"f1",  x"01",  x"7b", -- 02D8
         x"f1",  x"21",  x"7e",  x"f1",  x"cd",  x"6d",  x"12",  x"21", -- 02E0
         x"ae",  x"16",  x"22",  x"15",  x"f1",  x"3e",  x"45",  x"32", -- 02E8
         x"a6",  x"f1",  x"3e",  x"01",  x"32",  x"f5",  x"f0",  x"c9", -- 02F0
         x"2a",  x"08",  x"f1",  x"7e",  x"fe",  x"2f",  x"c2",  x"14", -- 02F8
         x"23",  x"3a",  x"9b",  x"f1",  x"b7",  x"c2",  x"0e",  x"23", -- 0300
         x"21",  x"5f",  x"17",  x"c3",  x"11",  x"23",  x"21",  x"3d", -- 0308
         x"17",  x"22",  x"08",  x"f1",  x"11",  x"6f",  x"f1",  x"cd", -- 0310
         x"37",  x"23",  x"23",  x"11",  x"5f",  x"f1",  x"cd",  x"37", -- 0318
         x"23",  x"23",  x"7e",  x"32",  x"f6",  x"f0",  x"23",  x"11", -- 0320
         x"83",  x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"08",  x"f1", -- 0328
         x"3a",  x"83",  x"f1",  x"32",  x"84",  x"f1",  x"c9",  x"06", -- 0330
         x"08",  x"1a",  x"86",  x"12",  x"13",  x"05",  x"c8",  x"78", -- 0338
         x"fe",  x"06",  x"c2",  x"39",  x"23",  x"13",  x"13",  x"c3", -- 0340
         x"39",  x"23",  x"3e",  x"01",  x"32",  x"0e",  x"f1",  x"3a", -- 0348
         x"9b",  x"f1",  x"b7",  x"c2",  x"65",  x"23",  x"06",  x"04", -- 0350
         x"21",  x"6b",  x"f1",  x"3a",  x"9d",  x"f1",  x"86",  x"77", -- 0358
         x"23",  x"05",  x"c2",  x"5b",  x"23",  x"0e",  x"02",  x"21", -- 0360
         x"77",  x"f1",  x"3a",  x"9d",  x"f1",  x"86",  x"77",  x"23", -- 0368
         x"0d",  x"c2",  x"6a",  x"23",  x"c9",  x"3e",  x"01",  x"32", -- 0370
         x"0e",  x"f1",  x"06",  x"02",  x"21",  x"61",  x"f1",  x"34", -- 0378
         x"23",  x"05",  x"c2",  x"7f",  x"23",  x"c9",  x"3e",  x"01", -- 0380
         x"32",  x"0f",  x"f1",  x"06",  x"02",  x"21",  x"5f",  x"f1", -- 0388
         x"34",  x"34",  x"23",  x"05",  x"c2",  x"90",  x"23",  x"c9", -- 0390
         x"2a",  x"a7",  x"f1",  x"7e",  x"fe",  x"2e",  x"c2",  x"ae", -- 0398
         x"23",  x"3a",  x"0b",  x"f1",  x"fe",  x"3b",  x"ca",  x"26", -- 03A0
         x"24",  x"af",  x"32",  x"82",  x"f1",  x"c9",  x"fe",  x"2f", -- 03A8
         x"c2",  x"c7",  x"23",  x"3a",  x"0b",  x"f1",  x"fe",  x"35", -- 03B0
         x"c2",  x"c1",  x"23",  x"21",  x"f2",  x"16",  x"c3",  x"c4", -- 03B8
         x"23",  x"21",  x"23",  x"17",  x"22",  x"a7",  x"f1",  x"3a", -- 03C0
         x"72",  x"f1",  x"86",  x"32",  x"72",  x"f1",  x"4e",  x"23", -- 03C8
         x"3a",  x"0b",  x"f1",  x"fe",  x"3b",  x"ca",  x"ed",  x"23", -- 03D0
         x"3a",  x"0e",  x"f1",  x"b7",  x"c2",  x"ed",  x"23",  x"3a", -- 03D8
         x"63",  x"f1",  x"86",  x"32",  x"63",  x"f1",  x"3a",  x"73", -- 03E0
         x"f1",  x"81",  x"32",  x"73",  x"f1",  x"3a",  x"62",  x"f1", -- 03E8
         x"86",  x"32",  x"62",  x"f1",  x"23",  x"7e",  x"32",  x"0f", -- 03F0
         x"f1",  x"23",  x"11",  x"82",  x"f1",  x"cd",  x"4d",  x"1b", -- 03F8
         x"22",  x"a7",  x"f1",  x"7e",  x"fe",  x"cc",  x"c0",  x"23", -- 0400
         x"22",  x"a7",  x"f1",  x"3a",  x"72",  x"f1",  x"c6",  x"0f", -- 0408
         x"32",  x"73",  x"f1",  x"3a",  x"62",  x"f1",  x"c6",  x"03", -- 0410
         x"32",  x"63",  x"f1",  x"3e",  x"44",  x"32",  x"83",  x"f1", -- 0418
         x"3e",  x"01",  x"32",  x"0e",  x"f1",  x"c9",  x"3e",  x"01", -- 0420
         x"32",  x"f6",  x"f0",  x"c9",  x"3e",  x"01",  x"32",  x"ec", -- 0428
         x"f0",  x"3a",  x"a3",  x"f0",  x"3d",  x"32",  x"a3",  x"f0", -- 0430
         x"f8",  x"32",  x"a7",  x"f0",  x"c9",  x"00",  x"3e",  x"0c", -- 0438
         x"32",  x"0b",  x"f1",  x"af",  x"32",  x"a6",  x"f1",  x"32", -- 0440
         x"14",  x"f1",  x"32",  x"1a",  x"f1",  x"32",  x"f8",  x"f0", -- 0448
         x"32",  x"f5",  x"f0",  x"32",  x"0a",  x"f1",  x"32",  x"eb", -- 0450
         x"f0",  x"32",  x"e9",  x"f0",  x"32",  x"ea",  x"f0",  x"32", -- 0458
         x"f1",  x"f0",  x"32",  x"00",  x"f1",  x"32",  x"f4",  x"f0", -- 0460
         x"32",  x"f3",  x"f0",  x"cd",  x"8c",  x"1a",  x"3e",  x"40", -- 0468
         x"32",  x"0e",  x"f1",  x"32",  x"ec",  x"f0",  x"3e",  x"01", -- 0470
         x"32",  x"19",  x"f1",  x"32",  x"e8",  x"f0",  x"3e",  x"09", -- 0478
         x"32",  x"f6",  x"f0",  x"32",  x"f7",  x"f0",  x"21",  x"84", -- 0480
         x"16",  x"22",  x"17",  x"f1",  x"21",  x"f2",  x"16",  x"22", -- 0488
         x"03",  x"f1",  x"3e",  x"fe",  x"32",  x"11",  x"f1",  x"3e", -- 0490
         x"02",  x"32",  x"12",  x"f1",  x"3e",  x"fd",  x"32",  x"1e", -- 0498
         x"f0",  x"3e",  x"bf",  x"32",  x"27",  x"f0",  x"32",  x"21", -- 04A0
         x"f0",  x"3e",  x"a7",  x"32",  x"24",  x"f0",  x"21",  x"e0", -- 04A8
         x"17",  x"22",  x"01",  x"f1",  x"01",  x"5b",  x"f1",  x"21", -- 04B0
         x"8a",  x"f1",  x"af",  x"cd",  x"6d",  x"12",  x"21",  x"bf", -- 04B8
         x"bf",  x"22",  x"5b",  x"f1",  x"21",  x"4f",  x"4f",  x"22", -- 04C0
         x"5d",  x"f1",  x"21",  x"a7",  x"a7",  x"22",  x"5f",  x"f1", -- 04C8
         x"21",  x"b7",  x"b7",  x"22",  x"61",  x"f1",  x"21",  x"6f", -- 04D0
         x"6f",  x"22",  x"63",  x"f1",  x"21",  x"7f",  x"7f",  x"22", -- 04D8
         x"65",  x"f1",  x"21",  x"67",  x"f1",  x"3e",  x"47",  x"77", -- 04E0
         x"23",  x"af",  x"77",  x"23",  x"3e",  x"47",  x"77",  x"23", -- 04E8
         x"af",  x"77",  x"23",  x"21",  x"5f",  x"6f",  x"22",  x"6b", -- 04F0
         x"f1",  x"21",  x"d7",  x"e7",  x"22",  x"6d",  x"f1",  x"21", -- 04F8
         x"00",  x"10",  x"22",  x"6f",  x"f1",  x"22",  x"71",  x"f1", -- 0500
         x"21",  x"a5",  x"b5",  x"22",  x"73",  x"f1",  x"22",  x"75", -- 0508
         x"f1",  x"21",  x"77",  x"f1",  x"3e",  x"c7",  x"77",  x"23", -- 0510
         x"af",  x"77",  x"23",  x"3e",  x"c7",  x"77",  x"23",  x"af", -- 0518
         x"77",  x"3e",  x"52",  x"57",  x"32",  x"fc",  x"f0",  x"cd", -- 0520
         x"66",  x"1a",  x"11",  x"7b",  x"f1",  x"cd",  x"82",  x"1a", -- 0528
         x"d5",  x"3e",  x"52",  x"57",  x"32",  x"fd",  x"f0",  x"cd", -- 0530
         x"66",  x"1a",  x"d1",  x"cd",  x"82",  x"1a",  x"d5",  x"3e", -- 0538
         x"46",  x"57",  x"32",  x"fa",  x"f0",  x"cd",  x"66",  x"1a", -- 0540
         x"d1",  x"cd",  x"82",  x"1a",  x"d5",  x"3e",  x"19",  x"57", -- 0548
         x"32",  x"fe",  x"f0",  x"cd",  x"66",  x"1a",  x"d1",  x"cd", -- 0550
         x"82",  x"1a",  x"af",  x"12",  x"32",  x"00",  x"f1",  x"13", -- 0558
         x"12",  x"32",  x"f4",  x"f0",  x"13",  x"d5",  x"3e",  x"11", -- 0560
         x"57",  x"32",  x"ff",  x"f0",  x"cd",  x"66",  x"1a",  x"d1", -- 0568
         x"cd",  x"82",  x"1a",  x"af",  x"12",  x"01",  x"8b",  x"f1", -- 0570
         x"21",  x"9a",  x"f1",  x"3e",  x"05",  x"cd",  x"6d",  x"12", -- 0578
         x"cd",  x"2a",  x"2c",  x"cd",  x"c0",  x"1d",  x"3a",  x"0b", -- 0580
         x"f1",  x"fe",  x"0c",  x"ca",  x"94",  x"25",  x"cd",  x"6f", -- 0588
         x"1b",  x"c3",  x"a0",  x"25",  x"cd",  x"3f",  x"1f",  x"cd", -- 0590
         x"82",  x"1b",  x"cd",  x"29",  x"2a",  x"cd",  x"b6",  x"2a", -- 0598
         x"cd",  x"eb",  x"28",  x"cd",  x"a9",  x"25",  x"c3",  x"80", -- 05A0
         x"25",  x"3a",  x"f5",  x"f0",  x"fe",  x"00",  x"ca",  x"b5", -- 05A8
         x"25",  x"3d",  x"32",  x"f5",  x"f0",  x"cd",  x"b6",  x"20", -- 05B0
         x"ca",  x"fa",  x"25",  x"32",  x"14",  x"f1",  x"47",  x"3a", -- 05B8
         x"a6",  x"f1",  x"fe",  x"00",  x"c2",  x"b7",  x"27",  x"32", -- 05C0
         x"14",  x"f1",  x"78",  x"32",  x"a6",  x"f1",  x"fe",  x"47", -- 05C8
         x"ca",  x"ef",  x"25",  x"fe",  x"4a",  x"ca",  x"12",  x"27", -- 05D0
         x"fe",  x"4c",  x"ca",  x"35",  x"27",  x"fe",  x"42",  x"ca", -- 05D8
         x"02",  x"27",  x"fe",  x"59",  x"ca",  x"1c",  x"27",  x"fe", -- 05E0
         x"53",  x"ca",  x"45",  x"27",  x"c3",  x"fa",  x"25",  x"3e", -- 05E8
         x"01",  x"32",  x"19",  x"f1",  x"21",  x"ac",  x"15",  x"c3", -- 05F0
         x"09",  x"26",  x"3a",  x"a6",  x"f1",  x"fe",  x"00",  x"c8", -- 05F8
         x"3a",  x"f5",  x"f0",  x"fe",  x"00",  x"c0",  x"2a",  x"15", -- 0600
         x"f1",  x"7e",  x"fe",  x"2f",  x"ca",  x"60",  x"26",  x"fe", -- 0608
         x"2e",  x"ca",  x"a2",  x"26",  x"11",  x"6f",  x"f1",  x"cd", -- 0610
         x"60",  x"1b",  x"23",  x"7e",  x"11",  x"5f",  x"f1",  x"cd", -- 0618
         x"60",  x"1b",  x"23",  x"7e",  x"32",  x"f5",  x"f0",  x"23", -- 0620
         x"11",  x"7f",  x"f1",  x"cd",  x"4d",  x"1b",  x"3a",  x"f9", -- 0628
         x"f0",  x"32",  x"fa",  x"f0",  x"22",  x"15",  x"f1",  x"7e", -- 0630
         x"fe",  x"cc",  x"c0",  x"23",  x"3a",  x"71",  x"f1",  x"86", -- 0638
         x"32",  x"7a",  x"f1",  x"23",  x"3a",  x"61",  x"f1",  x"86", -- 0640
         x"32",  x"6a",  x"f1",  x"23",  x"7e",  x"32",  x"f8",  x"f0", -- 0648
         x"3e",  x"05",  x"32",  x"9a",  x"f1",  x"23",  x"11",  x"8a", -- 0650
         x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"15",  x"f1",  x"c9", -- 0658
         x"3a",  x"a6",  x"f1",  x"fe",  x"52",  x"c2",  x"6e",  x"26", -- 0660
         x"21",  x"2a",  x"f0",  x"c3",  x"7b",  x"26",  x"fe",  x"54", -- 0668
         x"ca",  x"78",  x"26",  x"fe",  x"47",  x"c2",  x"81",  x"26", -- 0670
         x"21",  x"b0",  x"15",  x"22",  x"15",  x"f1",  x"c3",  x"09", -- 0678
         x"26",  x"fe",  x"46",  x"c2",  x"72",  x"1a",  x"21",  x"ce", -- 0680
         x"16",  x"c3",  x"7b",  x"26",  x"3e",  x"01",  x"32",  x"19", -- 0688
         x"f1",  x"32",  x"f5",  x"f0",  x"21",  x"2a",  x"f0",  x"22", -- 0690
         x"15",  x"f1",  x"3a",  x"14",  x"f1",  x"b7",  x"c8",  x"c3", -- 0698
         x"be",  x"25",  x"3a",  x"a6",  x"f1",  x"fe",  x"57",  x"ca", -- 06A0
         x"e7",  x"26",  x"fe",  x"46",  x"ca",  x"e7",  x"26",  x"fe", -- 06A8
         x"45",  x"ca",  x"e7",  x"26",  x"fe",  x"52",  x"ca",  x"8c", -- 06B0
         x"26",  x"fe",  x"59",  x"c2",  x"cc",  x"26",  x"3a",  x"ed", -- 06B8
         x"f0",  x"b7",  x"ca",  x"cc",  x"26",  x"af",  x"32",  x"ed", -- 06C0
         x"f0",  x"cd",  x"13",  x"f0",  x"af",  x"32",  x"a6",  x"f1", -- 06C8
         x"cd",  x"e3",  x"0f",  x"3e",  x"01",  x"32",  x"19",  x"f1", -- 06D0
         x"3a",  x"14",  x"f1",  x"47",  x"fe",  x"00",  x"c8",  x"af", -- 06D8
         x"32",  x"14",  x"f1",  x"78",  x"c3",  x"cb",  x"25",  x"cd", -- 06E0
         x"2c",  x"24",  x"af",  x"32",  x"a6",  x"f1",  x"cd",  x"e3", -- 06E8
         x"0f",  x"3a",  x"0b",  x"f1",  x"fe",  x"0a",  x"ca",  x"43", -- 06F0
         x"2c",  x"fe",  x"08",  x"ca",  x"fc",  x"2c",  x"cd",  x"56", -- 06F8
         x"20",  x"c9",  x"3a",  x"6f",  x"f1",  x"fe",  x"04",  x"d8", -- 0700
         x"af",  x"32",  x"19",  x"f1",  x"21",  x"e1",  x"15",  x"c3", -- 0708
         x"09",  x"26",  x"af",  x"32",  x"19",  x"f1",  x"21",  x"ef", -- 0710
         x"15",  x"c3",  x"09",  x"26",  x"af",  x"32",  x"19",  x"f1", -- 0718
         x"32",  x"ed",  x"f0",  x"3a",  x"fa",  x"f0",  x"fe",  x"3b", -- 0720
         x"3e",  x"fd",  x"ca",  x"2f",  x"27",  x"3e",  x"f8",  x"21", -- 0728
         x"c6",  x"15",  x"c3",  x"0a",  x"26",  x"3a",  x"fa",  x"f0", -- 0730
         x"fe",  x"3b",  x"c8",  x"af",  x"32",  x"19",  x"f1",  x"21", -- 0738
         x"7e",  x"16",  x"c3",  x"09",  x"26",  x"3a",  x"fa",  x"f0", -- 0740
         x"fe",  x"34",  x"ca",  x"52",  x"27",  x"fe",  x"36",  x"c2", -- 0748
         x"57",  x"27",  x"3e",  x"01",  x"c3",  x"77",  x"27",  x"fe", -- 0750
         x"3b",  x"c2",  x"66",  x"27",  x"3e",  x"05",  x"c3",  x"77", -- 0758
         x"27",  x"3e",  x"00",  x"c3",  x"77",  x"27",  x"fe",  x"35", -- 0760
         x"c2",  x"70",  x"27",  x"3e",  x"03",  x"c3",  x"77",  x"27", -- 0768
         x"fe",  x"37",  x"c2",  x"61",  x"27",  x"3e",  x"02",  x"11", -- 0770
         x"6f",  x"f1",  x"cd",  x"60",  x"1b",  x"32",  x"e7",  x"f0", -- 0778
         x"3a",  x"fa",  x"f0",  x"21",  x"ea",  x"16",  x"fe",  x"3b", -- 0780
         x"ca",  x"93",  x"27",  x"fe",  x"46",  x"ca",  x"93",  x"27", -- 0788
         x"21",  x"e6",  x"16",  x"3a",  x"e7",  x"f0",  x"11",  x"5f", -- 0790
         x"f1",  x"7e",  x"cd",  x"60",  x"1b",  x"23",  x"7e",  x"32", -- 0798
         x"f5",  x"f0",  x"23",  x"11",  x"7f",  x"f1",  x"cd",  x"4d", -- 07A0
         x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"fa",  x"f0",  x"22", -- 07A8
         x"15",  x"f1",  x"af",  x"32",  x"19",  x"f1",  x"c9",  x"3a", -- 07B0
         x"19",  x"f1",  x"b7",  x"ca",  x"fa",  x"25",  x"3a",  x"14", -- 07B8
         x"f1",  x"47",  x"af",  x"32",  x"14",  x"f1",  x"3a",  x"a6", -- 07C0
         x"f1",  x"fe",  x"52",  x"78",  x"c2",  x"0c",  x"28",  x"fe", -- 07C8
         x"53",  x"ca",  x"45",  x"27",  x"fe",  x"59",  x"ca",  x"1c", -- 07D0
         x"27",  x"fe",  x"4c",  x"ca",  x"35",  x"27",  x"fe",  x"42", -- 07D8
         x"ca",  x"fa",  x"25",  x"fe",  x"47",  x"ca",  x"ed",  x"27", -- 07E0
         x"fe",  x"4a",  x"c2",  x"0c",  x"28",  x"3a",  x"e8",  x"f0", -- 07E8
         x"b7",  x"ca",  x"fa",  x"25",  x"3a",  x"1a",  x"f1",  x"b7", -- 07F0
         x"3a",  x"e8",  x"f0",  x"ca",  x"06",  x"28",  x"fe",  x"01", -- 07F8
         x"ca",  x"0b",  x"28",  x"c3",  x"fa",  x"25",  x"fe",  x"01", -- 0800
         x"ca",  x"fa",  x"25",  x"78",  x"32",  x"a6",  x"f1",  x"fe", -- 0808
         x"4c",  x"ca",  x"91",  x"28",  x"fe",  x"4a",  x"ca",  x"1e", -- 0810
         x"28",  x"fe",  x"59",  x"c2",  x"ce",  x"25",  x"3a",  x"fa", -- 0818
         x"f0",  x"fe",  x"46",  x"ca",  x"ca",  x"25",  x"fe",  x"36", -- 0820
         x"ca",  x"30",  x"28",  x"fe",  x"34",  x"c2",  x"73",  x"28", -- 0828
         x"3e",  x"01",  x"11",  x"6f",  x"f1",  x"cd",  x"60",  x"1b", -- 0830
         x"af",  x"32",  x"19",  x"f1",  x"3e",  x"00",  x"11",  x"5f", -- 0838
         x"f1",  x"cd",  x"60",  x"1b",  x"3e",  x"07",  x"32",  x"f5", -- 0840
         x"f0",  x"21",  x"c1",  x"15",  x"3a",  x"a6",  x"f1",  x"fe", -- 0848
         x"59",  x"ca",  x"57",  x"28",  x"21",  x"ea",  x"15",  x"11", -- 0850
         x"7f",  x"f1",  x"3a",  x"fa",  x"f0",  x"fe",  x"3b",  x"c2", -- 0858
         x"66",  x"28",  x"01",  x"04",  x"00",  x"09",  x"cd",  x"4d", -- 0860
         x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"fa",  x"f0",  x"22", -- 0868
         x"15",  x"f1",  x"c9",  x"fe",  x"3b",  x"c2",  x"7d",  x"28", -- 0870
         x"3e",  x"05",  x"c3",  x"32",  x"28",  x"fe",  x"35",  x"c2", -- 0878
         x"87",  x"28",  x"3e",  x"03",  x"c3",  x"32",  x"28",  x"fe", -- 0880
         x"37",  x"c2",  x"30",  x"28",  x"3e",  x"02",  x"c3",  x"32", -- 0888
         x"28",  x"3a",  x"fa",  x"f0",  x"fe",  x"34",  x"ca",  x"9e", -- 0890
         x"28",  x"fe",  x"36",  x"c2",  x"ca",  x"28",  x"3e",  x"fc", -- 0898
         x"11",  x"6f",  x"f1",  x"cd",  x"60",  x"1b",  x"af",  x"32", -- 08A0
         x"19",  x"f1",  x"3e",  x"00",  x"11",  x"5f",  x"f1",  x"cd", -- 08A8
         x"60",  x"1b",  x"3e",  x"0b",  x"32",  x"f5",  x"f0",  x"21", -- 08B0
         x"81",  x"16",  x"11",  x"7f",  x"f1",  x"cd",  x"4d",  x"1b", -- 08B8
         x"3a",  x"f9",  x"f0",  x"32",  x"fa",  x"f0",  x"22",  x"15", -- 08C0
         x"f1",  x"c9",  x"fe",  x"35",  x"ca",  x"d4",  x"28",  x"fe", -- 08C8
         x"37",  x"c2",  x"d9",  x"28",  x"3e",  x"00",  x"c3",  x"a0", -- 08D0
         x"28",  x"fe",  x"46",  x"c2",  x"e3",  x"28",  x"3e",  x"fb", -- 08D8
         x"c3",  x"a0",  x"28",  x"fe",  x"3b",  x"c2",  x"45",  x"27", -- 08E0
         x"c3",  x"fa",  x"25",  x"3a",  x"fe",  x"f0",  x"b7",  x"ca", -- 08E8
         x"6b",  x"29",  x"3a",  x"ea",  x"f0",  x"b7",  x"c2",  x"16", -- 08F0
         x"29",  x"3a",  x"f4",  x"f0",  x"b7",  x"c2",  x"16",  x"29", -- 08F8
         x"3a",  x"05",  x"f1",  x"b7",  x"ca",  x"0e",  x"29",  x"3d", -- 0900
         x"32",  x"05",  x"f1",  x"c2",  x"16",  x"29",  x"3e",  x"01", -- 0908
         x"32",  x"e9",  x"f0",  x"cd",  x"8c",  x"1a",  x"3a",  x"f6", -- 0910
         x"f0",  x"fe",  x"00",  x"ca",  x"27",  x"29",  x"3d",  x"32", -- 0918
         x"f6",  x"f0",  x"fe",  x"00",  x"c2",  x"6b",  x"29",  x"2a", -- 0920
         x"17",  x"f1",  x"7e",  x"fe",  x"2f",  x"c2",  x"36",  x"29", -- 0928
         x"21",  x"84",  x"16",  x"c3",  x"2a",  x"29",  x"fe",  x"2e", -- 0930
         x"c2",  x"48",  x"29",  x"af",  x"32",  x"ea",  x"f0",  x"32", -- 0938
         x"83",  x"f1",  x"32",  x"fe",  x"f0",  x"c3",  x"6b",  x"29", -- 0940
         x"11",  x"73",  x"f1",  x"cd",  x"60",  x"1b",  x"23",  x"7e", -- 0948
         x"11",  x"63",  x"f1",  x"cd",  x"60",  x"1b",  x"23",  x"7e", -- 0950
         x"32",  x"f6",  x"f0",  x"23",  x"11",  x"83",  x"f1",  x"cd", -- 0958
         x"4d",  x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"fe",  x"f0", -- 0960
         x"22",  x"17",  x"f1",  x"3a",  x"f3",  x"f0",  x"b7",  x"ca", -- 0968
         x"ab",  x"29",  x"3d",  x"32",  x"f3",  x"f0",  x"b7",  x"c0", -- 0970
         x"3a",  x"f4",  x"f0",  x"fe",  x"27",  x"c2",  x"81",  x"29", -- 0978
         x"c9",  x"2a",  x"08",  x"f1",  x"7e",  x"fe",  x"2f",  x"c2", -- 0980
         x"8d",  x"29",  x"21",  x"e2",  x"16",  x"3a",  x"78",  x"f1", -- 0988
         x"cd",  x"1a",  x"f0",  x"32",  x"78",  x"f1",  x"3e",  x"01", -- 0990
         x"32",  x"f3",  x"f0",  x"11",  x"88",  x"f1",  x"cd",  x"4d", -- 0998
         x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"f4",  x"f0",  x"22", -- 09A0
         x"08",  x"f1",  x"c9",  x"3a",  x"e9",  x"f0",  x"b7",  x"c8", -- 09A8
         x"3a",  x"ea",  x"f0",  x"b7",  x"c0",  x"3a",  x"fe",  x"f0", -- 09B0
         x"b7",  x"c8",  x"3a",  x"f4",  x"f0",  x"b7",  x"c0",  x"3a", -- 09B8
         x"fe",  x"f0",  x"fe",  x"1d",  x"ca",  x"ca",  x"29",  x"fe", -- 09C0
         x"4e",  x"c0",  x"3a",  x"0b",  x"f1",  x"fe",  x"0c",  x"c2", -- 09C8
         x"1a",  x"2a",  x"3a",  x"a4",  x"f0",  x"b7",  x"e2",  x"1a", -- 09D0
         x"2a",  x"3e",  x"09",  x"32",  x"98",  x"f1",  x"3e",  x"02", -- 09D8
         x"32",  x"1b",  x"f0",  x"06",  x"08",  x"3a",  x"73",  x"f1", -- 09E0
         x"80",  x"32",  x"78",  x"f1",  x"3a",  x"0a",  x"f1",  x"b7", -- 09E8
         x"06",  x"10",  x"3a",  x"63",  x"f1",  x"e2",  x"fa",  x"29", -- 09F0
         x"06",  x"08",  x"80",  x"32",  x"68",  x"f1",  x"11",  x"88", -- 09F8
         x"f1",  x"21",  x"e2",  x"16",  x"cd",  x"4d",  x"1b",  x"3a", -- 0A00
         x"f9",  x"f0",  x"32",  x"f4",  x"f0",  x"22",  x"08",  x"f1", -- 0A08
         x"3e",  x"01",  x"32",  x"f3",  x"f0",  x"af",  x"32",  x"e9", -- 0A10
         x"f0",  x"c9",  x"3e",  x"05",  x"32",  x"98",  x"f1",  x"3e", -- 0A18
         x"fe",  x"32",  x"1b",  x"f0",  x"06",  x"00",  x"c3",  x"e5", -- 0A20
         x"29",  x"3a",  x"0e",  x"f1",  x"fe",  x"00",  x"ca",  x"36", -- 0A28
         x"2a",  x"3d",  x"32",  x"0e",  x"f1",  x"c0",  x"3a",  x"5b", -- 0A30
         x"f1",  x"47",  x"3a",  x"11",  x"f1",  x"80",  x"32",  x"5b", -- 0A38
         x"f1",  x"32",  x"5c",  x"f1",  x"3a",  x"5d",  x"f1",  x"47", -- 0A40
         x"3a",  x"12",  x"f1",  x"80",  x"32",  x"5d",  x"f1",  x"32", -- 0A48
         x"5e",  x"f1",  x"3a",  x"a6",  x"f1",  x"fe",  x"54",  x"ca", -- 0A50
         x"5f",  x"2a",  x"fe",  x"52",  x"c2",  x"7b",  x"2a",  x"3a", -- 0A58
         x"1a",  x"f1",  x"b7",  x"3a",  x"11",  x"f1",  x"ca",  x"6c", -- 0A60
         x"2a",  x"3a",  x"12",  x"f1",  x"47",  x"3a",  x"6a",  x"f1", -- 0A68
         x"80",  x"32",  x"6a",  x"f1",  x"78",  x"11",  x"5f",  x"f1", -- 0A70
         x"cd",  x"60",  x"1b",  x"3a",  x"5d",  x"f1",  x"fe",  x"4f", -- 0A78
         x"ca",  x"88",  x"2a",  x"fe",  x"bf",  x"c2",  x"9b",  x"2a", -- 0A80
         x"3a",  x"11",  x"f1",  x"2f",  x"3c",  x"32",  x"11",  x"f1", -- 0A88
         x"3a",  x"12",  x"f1",  x"2f",  x"3c",  x"32",  x"12",  x"f1", -- 0A90
         x"c3",  x"a2",  x"2a",  x"fe",  x"87",  x"3e",  x"01",  x"c2", -- 0A98
         x"a8",  x"2a",  x"3e",  x"40",  x"32",  x"0e",  x"f1",  x"c9", -- 0AA0
         x"32",  x"0e",  x"f1",  x"3a",  x"a6",  x"f1",  x"fe",  x"52", -- 0AA8
         x"c0",  x"af",  x"32",  x"e8",  x"f0",  x"c9",  x"3a",  x"ff", -- 0AB0
         x"f0",  x"b7",  x"c8",  x"3a",  x"f1",  x"f0",  x"b7",  x"c2", -- 0AB8
         x"40",  x"2b",  x"3a",  x"eb",  x"f0",  x"b7",  x"c2",  x"e9", -- 0AC0
         x"2a",  x"2a",  x"01",  x"f1",  x"3a",  x"0a",  x"f1",  x"be", -- 0AC8
         x"c2",  x"40",  x"2b",  x"3e",  x"01",  x"32",  x"eb",  x"f0", -- 0AD0
         x"23",  x"7e",  x"fe",  x"ff",  x"c2",  x"e2",  x"2a",  x"21", -- 0AD8
         x"e0",  x"17",  x"22",  x"01",  x"f1",  x"af",  x"32",  x"0a", -- 0AE0
         x"f1",  x"3a",  x"00",  x"f1",  x"b7",  x"c2",  x"40",  x"2b", -- 0AE8
         x"3a",  x"ff",  x"f0",  x"fe",  x"14",  x"06",  x"08",  x"c2", -- 0AF0
         x"40",  x"2b",  x"3a",  x"99",  x"f1",  x"fe",  x"05",  x"78", -- 0AF8
         x"ca",  x"05",  x"2b",  x"2f",  x"3c",  x"47",  x"3a",  x"79", -- 0B00
         x"f1",  x"80",  x"47",  x"fe",  x"7d",  x"d2",  x"15",  x"2b", -- 0B08
         x"3e",  x"09",  x"c3",  x"1c",  x"2b",  x"fe",  x"c8",  x"da", -- 0B10
         x"25",  x"2b",  x"3e",  x"05",  x"32",  x"99",  x"f1",  x"32", -- 0B18
         x"97",  x"f1",  x"c3",  x"28",  x"2b",  x"32",  x"79",  x"f1", -- 0B20
         x"3e",  x"0a",  x"32",  x"f7",  x"f0",  x"21",  x"13",  x"17", -- 0B28
         x"11",  x"89",  x"f1",  x"cd",  x"4d",  x"1b",  x"3a",  x"f9", -- 0B30
         x"f0",  x"32",  x"ff",  x"f0",  x"22",  x"03",  x"f1",  x"c9", -- 0B38
         x"3a",  x"f7",  x"f0",  x"fe",  x"00",  x"c2",  x"50",  x"2b", -- 0B40
         x"3a",  x"eb",  x"f0",  x"b7",  x"c8",  x"c3",  x"57",  x"2b", -- 0B48
         x"3d",  x"32",  x"f7",  x"f0",  x"fe",  x"00",  x"c0",  x"2a", -- 0B50
         x"03",  x"f1",  x"7e",  x"fe",  x"2f",  x"c2",  x"66",  x"2b", -- 0B58
         x"21",  x"f2",  x"16",  x"c3",  x"5a",  x"2b",  x"fe",  x"2e", -- 0B60
         x"ca",  x"03",  x"2c",  x"3a",  x"99",  x"f1",  x"fe",  x"05", -- 0B68
         x"7e",  x"ca",  x"76",  x"2b",  x"2f",  x"3c",  x"47",  x"3a", -- 0B70
         x"79",  x"f1",  x"80",  x"47",  x"23",  x"3a",  x"69",  x"f1", -- 0B78
         x"86",  x"32",  x"69",  x"f1",  x"23",  x"7e",  x"32",  x"f7", -- 0B80
         x"f0",  x"23",  x"11",  x"89",  x"f1",  x"cd",  x"4d",  x"1b", -- 0B88
         x"3a",  x"f9",  x"f0",  x"32",  x"ff",  x"f0",  x"22",  x"03", -- 0B90
         x"f1",  x"78",  x"fe",  x"7d",  x"d2",  x"a9",  x"2b",  x"3e", -- 0B98
         x"02",  x"32",  x"1e",  x"f0",  x"3e",  x"09",  x"c3",  x"b5", -- 0BA0
         x"2b",  x"fe",  x"c8",  x"da",  x"be",  x"2b",  x"3e",  x"fe", -- 0BA8
         x"32",  x"1e",  x"f0",  x"3e",  x"05",  x"32",  x"99",  x"f1", -- 0BB0
         x"32",  x"97",  x"f1",  x"c3",  x"c1",  x"2b",  x"32",  x"79", -- 0BB8
         x"f1",  x"3a",  x"79",  x"f1",  x"32",  x"77",  x"f1",  x"3a", -- 0BC0
         x"69",  x"f1",  x"32",  x"67",  x"f1",  x"7e",  x"fe",  x"cc", -- 0BC8
         x"c0",  x"23",  x"3a",  x"99",  x"f1",  x"fe",  x"05",  x"7e", -- 0BD0
         x"ca",  x"dd",  x"2b",  x"2f",  x"3c",  x"47",  x"3a",  x"77", -- 0BD8
         x"f1",  x"80",  x"32",  x"77",  x"f1",  x"23",  x"3a",  x"67", -- 0BE0
         x"f1",  x"86",  x"32",  x"67",  x"f1",  x"23",  x"7e",  x"32", -- 0BE8
         x"f7",  x"f0",  x"23",  x"11",  x"87",  x"f1",  x"cd",  x"4d", -- 0BF0
         x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"00",  x"f1",  x"22", -- 0BF8
         x"03",  x"f1",  x"c9",  x"3a",  x"f1",  x"f0",  x"b7",  x"ca", -- 0C00
         x"1b",  x"2c",  x"af",  x"32",  x"ff",  x"f0",  x"32",  x"89", -- 0C08
         x"f1",  x"32",  x"f1",  x"f0",  x"32",  x"eb",  x"f0",  x"32", -- 0C10
         x"f7",  x"f0",  x"c9",  x"3a",  x"77",  x"f1",  x"cd",  x"1d", -- 0C18
         x"f0",  x"32",  x"77",  x"f1",  x"3e",  x"01",  x"32",  x"f7", -- 0C20
         x"f0",  x"c9",  x"cd",  x"9f",  x"1a",  x"3a",  x"f8",  x"f0", -- 0C28
         x"fe",  x"00",  x"c8",  x"3d",  x"32",  x"f8",  x"f0",  x"c0", -- 0C30
         x"af",  x"32",  x"8a",  x"f1",  x"c9",  x"00",  x"3e",  x"0a", -- 0C38
         x"32",  x"0b",  x"f1",  x"af",  x"32",  x"a6",  x"f1",  x"32", -- 0C40
         x"14",  x"f1",  x"32",  x"f8",  x"f0",  x"32",  x"f5",  x"f0", -- 0C48
         x"32",  x"0a",  x"f1",  x"32",  x"eb",  x"f0",  x"32",  x"e9", -- 0C50
         x"f0",  x"32",  x"ea",  x"f0",  x"32",  x"f4",  x"f0",  x"32", -- 0C58
         x"f3",  x"f0",  x"cd",  x"8c",  x"1a",  x"3e",  x"01",  x"32", -- 0C60
         x"19",  x"f1",  x"32",  x"e8",  x"f0",  x"32",  x"ec",  x"f0", -- 0C68
         x"3e",  x"09",  x"32",  x"f6",  x"f0",  x"21",  x"84",  x"16", -- 0C70
         x"22",  x"17",  x"f1",  x"01",  x"5b",  x"f1",  x"21",  x"8a", -- 0C78
         x"f1",  x"af",  x"cd",  x"6d",  x"12",  x"21",  x"93",  x"93", -- 0C80
         x"22",  x"5f",  x"f1",  x"22",  x"63",  x"f1",  x"21",  x"a3", -- 0C88
         x"a3",  x"22",  x"61",  x"f1",  x"22",  x"65",  x"f1",  x"21", -- 0C90
         x"67",  x"f1",  x"af",  x"77",  x"23",  x"77",  x"21",  x"00", -- 0C98
         x"10",  x"22",  x"6f",  x"f1",  x"22",  x"71",  x"f1",  x"21", -- 0CA0
         x"c5",  x"d5",  x"22",  x"73",  x"f1",  x"22",  x"75",  x"f1", -- 0CA8
         x"21",  x"77",  x"f1",  x"af",  x"77",  x"23",  x"77",  x"3e", -- 0CB0
         x"46",  x"57",  x"32",  x"fa",  x"f0",  x"cd",  x"66",  x"1a", -- 0CB8
         x"11",  x"7f",  x"f1",  x"cd",  x"82",  x"1a",  x"d5",  x"3e", -- 0CC0
         x"19",  x"57",  x"32",  x"fe",  x"f0",  x"cd",  x"66",  x"1a", -- 0CC8
         x"d1",  x"cd",  x"82",  x"1a",  x"af",  x"12",  x"13",  x"12", -- 0CD0
         x"01",  x"8b",  x"f1",  x"21",  x"9a",  x"f1",  x"3e",  x"05", -- 0CD8
         x"cd",  x"6d",  x"12",  x"c3",  x"80",  x"25",  x"00",  x"cd", -- 0CE0
         x"77",  x"14",  x"3e",  x"08",  x"32",  x"0b",  x"f1",  x"32", -- 0CE8
         x"ec",  x"f0",  x"af",  x"01",  x"5b",  x"f1",  x"21",  x"8a", -- 0CF0
         x"f1",  x"cd",  x"6d",  x"12",  x"af",  x"32",  x"a6",  x"f1", -- 0CF8
         x"32",  x"14",  x"f1",  x"32",  x"f8",  x"f0",  x"32",  x"f5", -- 0D00
         x"f0",  x"32",  x"eb",  x"f0",  x"32",  x"fe",  x"f0",  x"3e", -- 0D08
         x"01",  x"32",  x"0e",  x"f1",  x"32",  x"19",  x"f1",  x"3c", -- 0D10
         x"32",  x"0f",  x"f1",  x"3c",  x"32",  x"10",  x"f1",  x"21", -- 0D18
         x"ae",  x"34",  x"22",  x"17",  x"f1",  x"22",  x"08",  x"f1", -- 0D20
         x"22",  x"03",  x"f1",  x"21",  x"e0",  x"17",  x"7e",  x"32", -- 0D28
         x"ee",  x"f0",  x"23",  x"7e",  x"32",  x"ef",  x"f0",  x"23", -- 0D30
         x"7e",  x"32",  x"f0",  x"f0",  x"22",  x"06",  x"f1",  x"21", -- 0D38
         x"92",  x"92",  x"22",  x"5f",  x"f1",  x"21",  x"a2",  x"a2", -- 0D40
         x"22",  x"61",  x"f1",  x"21",  x"ab",  x"ab",  x"22",  x"5b", -- 0D48
         x"f1",  x"22",  x"63",  x"f1",  x"22",  x"66",  x"f1",  x"3e", -- 0D50
         x"ab",  x"32",  x"5d",  x"f1",  x"32",  x"65",  x"f1",  x"32", -- 0D58
         x"68",  x"f1",  x"21",  x"00",  x"10",  x"22",  x"6f",  x"f1", -- 0D60
         x"22",  x"71",  x"f1",  x"21",  x"30",  x"40",  x"22",  x"6b", -- 0D68
         x"f1",  x"21",  x"60",  x"70",  x"22",  x"73",  x"f1",  x"21", -- 0D70
         x"90",  x"a0",  x"22",  x"76",  x"f1",  x"3e",  x"38",  x"32", -- 0D78
         x"6d",  x"f1",  x"3e",  x"68",  x"32",  x"75",  x"f1",  x"3e", -- 0D80
         x"98",  x"32",  x"78",  x"f1",  x"3e",  x"3e",  x"57",  x"cd", -- 0D88
         x"66",  x"1a",  x"11",  x"7b",  x"f1",  x"cd",  x"82",  x"1a", -- 0D90
         x"3e",  x"3e",  x"57",  x"cd",  x"66",  x"1a",  x"11",  x"83", -- 0D98
         x"f1",  x"cd",  x"82",  x"1a",  x"3e",  x"3e",  x"57",  x"cd", -- 0DA0
         x"66",  x"1a",  x"11",  x"86",  x"f1",  x"cd",  x"82",  x"1a", -- 0DA8
         x"3e",  x"46",  x"32",  x"fa",  x"f0",  x"57",  x"cd",  x"66", -- 0DB0
         x"1a",  x"11",  x"7f",  x"f1",  x"cd",  x"82",  x"1a",  x"01", -- 0DB8
         x"8b",  x"f1",  x"21",  x"9a",  x"f1",  x"3e",  x"05",  x"cd", -- 0DC0
         x"6d",  x"12",  x"cd",  x"2a",  x"2c",  x"cd",  x"91",  x"2f", -- 0DC8
         x"cd",  x"d9",  x"2d",  x"cd",  x"a9",  x"25",  x"c3",  x"ca", -- 0DD0
         x"2d",  x"3a",  x"0e",  x"f1",  x"3d",  x"32",  x"0e",  x"f1", -- 0DD8
         x"c2",  x"6c",  x"2e",  x"2a",  x"17",  x"f1",  x"7e",  x"fe", -- 0DE0
         x"2f",  x"c2",  x"52",  x"2e",  x"3a",  x"eb",  x"f0",  x"b7", -- 0DE8
         x"ca",  x"fe",  x"2d",  x"fe",  x"01",  x"c2",  x"fe",  x"2d", -- 0DF0
         x"21",  x"bc",  x"34",  x"c3",  x"52",  x"2e",  x"23",  x"22", -- 0DF8
         x"17",  x"f1",  x"3a",  x"ee",  x"f0",  x"3d",  x"32",  x"ee", -- 0E00
         x"f0",  x"11",  x"f3",  x"ff",  x"19",  x"c2",  x"52",  x"2e", -- 0E08
         x"2a",  x"06",  x"f1",  x"3a",  x"7d",  x"f1",  x"fe",  x"58", -- 0E10
         x"3e",  x"00",  x"c2",  x"1f",  x"2e",  x"3e",  x"10",  x"86", -- 0E18
         x"32",  x"ee",  x"f0",  x"23",  x"7e",  x"fe",  x"ff",  x"c2", -- 0E20
         x"2d",  x"2e",  x"21",  x"e0",  x"17",  x"22",  x"06",  x"f1", -- 0E28
         x"2a",  x"17",  x"f1",  x"7e",  x"fe",  x"2e",  x"ca",  x"44", -- 0E30
         x"2e",  x"3a",  x"5b",  x"f1",  x"c6",  x"08",  x"32",  x"5b", -- 0E38
         x"f1",  x"c3",  x"52",  x"2e",  x"3a",  x"5b",  x"f1",  x"c6", -- 0E40
         x"f0",  x"32",  x"5b",  x"f1",  x"32",  x"5c",  x"f1",  x"21", -- 0E48
         x"94",  x"34",  x"23",  x"3a",  x"5b",  x"f1",  x"86",  x"32", -- 0E50
         x"5b",  x"f1",  x"32",  x"5c",  x"f1",  x"23",  x"7e",  x"32", -- 0E58
         x"0e",  x"f1",  x"23",  x"11",  x"7b",  x"f1",  x"cd",  x"4d", -- 0E60
         x"1b",  x"22",  x"17",  x"f1",  x"3a",  x"0f",  x"f1",  x"3d", -- 0E68
         x"32",  x"0f",  x"f1",  x"c2",  x"ff",  x"2e",  x"2a",  x"08", -- 0E70
         x"f1",  x"7e",  x"fe",  x"2f",  x"c2",  x"e5",  x"2e",  x"3a", -- 0E78
         x"eb",  x"f0",  x"b7",  x"ca",  x"91",  x"2e",  x"fe",  x"02", -- 0E80
         x"c2",  x"91",  x"2e",  x"21",  x"bc",  x"34",  x"c3",  x"e5", -- 0E88
         x"2e",  x"23",  x"22",  x"08",  x"f1",  x"3a",  x"ef",  x"f0", -- 0E90
         x"3d",  x"32",  x"ef",  x"f0",  x"11",  x"f3",  x"ff",  x"19", -- 0E98
         x"c2",  x"e5",  x"2e",  x"2a",  x"06",  x"f1",  x"3a",  x"85", -- 0EA0
         x"f1",  x"fe",  x"58",  x"3e",  x"00",  x"c2",  x"b2",  x"2e", -- 0EA8
         x"3e",  x"10",  x"86",  x"32",  x"ef",  x"f0",  x"23",  x"7e", -- 0EB0
         x"fe",  x"ff",  x"c2",  x"c0",  x"2e",  x"21",  x"e0",  x"17", -- 0EB8
         x"22",  x"06",  x"f1",  x"2a",  x"08",  x"f1",  x"7e",  x"fe", -- 0EC0
         x"2e",  x"ca",  x"d7",  x"2e",  x"3a",  x"63",  x"f1",  x"c6", -- 0EC8
         x"08",  x"32",  x"63",  x"f1",  x"c3",  x"e5",  x"2e",  x"3a", -- 0ED0
         x"63",  x"f1",  x"c6",  x"f0",  x"32",  x"63",  x"f1",  x"32", -- 0ED8
         x"64",  x"f1",  x"21",  x"94",  x"34",  x"23",  x"3a",  x"63", -- 0EE0
         x"f1",  x"86",  x"32",  x"63",  x"f1",  x"32",  x"64",  x"f1", -- 0EE8
         x"23",  x"7e",  x"32",  x"0f",  x"f1",  x"23",  x"11",  x"83", -- 0EF0
         x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"08",  x"f1",  x"3a", -- 0EF8
         x"10",  x"f1",  x"3d",  x"32",  x"10",  x"f1",  x"c0",  x"2a", -- 0F00
         x"03",  x"f1",  x"7e",  x"fe",  x"2f",  x"c2",  x"76",  x"2f", -- 0F08
         x"3a",  x"eb",  x"f0",  x"b7",  x"ca",  x"22",  x"2f",  x"fe", -- 0F10
         x"03",  x"c2",  x"22",  x"2f",  x"21",  x"bc",  x"34",  x"c3", -- 0F18
         x"76",  x"2f",  x"23",  x"22",  x"03",  x"f1",  x"3a",  x"f0", -- 0F20
         x"f0",  x"3d",  x"32",  x"f0",  x"f0",  x"11",  x"f3",  x"ff", -- 0F28
         x"19",  x"c2",  x"76",  x"2f",  x"2a",  x"06",  x"f1",  x"3a", -- 0F30
         x"88",  x"f1",  x"fe",  x"58",  x"3e",  x"00",  x"c2",  x"43", -- 0F38
         x"2f",  x"3e",  x"10",  x"86",  x"32",  x"f0",  x"f0",  x"23", -- 0F40
         x"7e",  x"fe",  x"ff",  x"c2",  x"51",  x"2f",  x"21",  x"e0", -- 0F48
         x"17",  x"22",  x"06",  x"f1",  x"2a",  x"03",  x"f1",  x"7e", -- 0F50
         x"fe",  x"2e",  x"ca",  x"68",  x"2f",  x"3a",  x"66",  x"f1", -- 0F58
         x"c6",  x"08",  x"32",  x"66",  x"f1",  x"c3",  x"76",  x"2f", -- 0F60
         x"3a",  x"66",  x"f1",  x"c6",  x"f0",  x"32",  x"66",  x"f1", -- 0F68
         x"32",  x"67",  x"f1",  x"21",  x"94",  x"34",  x"23",  x"3a", -- 0F70
         x"66",  x"f1",  x"86",  x"32",  x"66",  x"f1",  x"32",  x"67", -- 0F78
         x"f1",  x"23",  x"7e",  x"32",  x"10",  x"f1",  x"23",  x"11", -- 0F80
         x"86",  x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"03",  x"f1", -- 0F88
         x"c9",  x"3a",  x"6f",  x"f1",  x"fe",  x"e0",  x"da",  x"a0", -- 0F90
         x"2f",  x"fe",  x"f0",  x"d2",  x"a0",  x"2f",  x"c1",  x"c9", -- 0F98
         x"3a",  x"a6",  x"f1",  x"fe",  x"57",  x"c8",  x"fe",  x"4a", -- 0FA0
         x"ca",  x"5c",  x"30",  x"3a",  x"eb",  x"f0",  x"b7",  x"ca", -- 0FA8
         x"db",  x"2f",  x"fe",  x"04",  x"ca",  x"db",  x"2f",  x"3a", -- 0FB0
         x"6f",  x"f1",  x"fe",  x"2a",  x"da",  x"e4",  x"2f",  x"fe", -- 0FB8
         x"3d",  x"d8",  x"fe",  x"5a",  x"da",  x"e4",  x"2f",  x"fe", -- 0FC0
         x"6d",  x"d8",  x"fe",  x"8a",  x"da",  x"e4",  x"2f",  x"fe", -- 0FC8
         x"9d",  x"d8",  x"fe",  x"a0",  x"d8",  x"fe",  x"b0",  x"da", -- 0FD0
         x"e4",  x"2f",  x"c9",  x"3a",  x"6f",  x"f1",  x"fe",  x"15", -- 0FD8
         x"d8",  x"fe",  x"ba",  x"d0",  x"af",  x"32",  x"19",  x"f1", -- 0FE0
         x"3e",  x"09",  x"32",  x"f5",  x"f0",  x"21",  x"a8",  x"a8", -- 0FE8
         x"22",  x"5f",  x"f1",  x"22",  x"61",  x"f1",  x"3a",  x"eb", -- 0FF0
         x"f0",  x"b7",  x"c2",  x"09",  x"30",  x"21",  x"20",  x"30", -- 0FF8
         x"22",  x"6f",  x"f1",  x"22",  x"71",  x"f1",  x"c3",  x"19", -- 1000
         x"30",  x"3a",  x"a6",  x"f1",  x"fe",  x"42",  x"c2",  x"19", -- 1008
         x"30",  x"3e",  x"f0",  x"11",  x"6f",  x"f1",  x"cd",  x"60", -- 1010
         x"1b",  x"3e",  x"57",  x"32",  x"a6",  x"f1",  x"3a",  x"eb", -- 1018
         x"f0",  x"fe",  x"04",  x"ca",  x"42",  x"30",  x"b7",  x"ca", -- 1020
         x"42",  x"30",  x"21",  x"a3",  x"a3",  x"22",  x"5b",  x"f1", -- 1028
         x"22",  x"63",  x"f1",  x"22",  x"66",  x"f1",  x"21",  x"a1", -- 1030
         x"34",  x"22",  x"17",  x"f1",  x"22",  x"08",  x"f1",  x"22", -- 1038
         x"03",  x"f1",  x"af",  x"32",  x"eb",  x"f0",  x"cd",  x"e3", -- 1040
         x"0f",  x"21",  x"9a",  x"15",  x"11",  x"7f",  x"f1",  x"cd", -- 1048
         x"4d",  x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"fa",  x"f0", -- 1050
         x"22",  x"15",  x"f1",  x"c9",  x"3a",  x"fa",  x"f0",  x"fe", -- 1058
         x"49",  x"c0",  x"3a",  x"eb",  x"f0",  x"fe",  x"04",  x"c8", -- 1060
         x"b7",  x"c2",  x"b3",  x"30",  x"3a",  x"6f",  x"f1",  x"fe", -- 1068
         x"18",  x"d2",  x"80",  x"30",  x"fe",  x"08",  x"d8",  x"3a", -- 1070
         x"5f",  x"f1",  x"fe",  x"90",  x"d8",  x"c3",  x"e4",  x"2f", -- 1078
         x"3a",  x"7d",  x"f1",  x"b7",  x"c2",  x"77",  x"30",  x"3a", -- 1080
         x"5f",  x"f1",  x"47",  x"3a",  x"5b",  x"f1",  x"90",  x"fe", -- 1088
         x"1f",  x"c0",  x"21",  x"8b",  x"8b",  x"22",  x"5f",  x"f1", -- 1090
         x"21",  x"9b",  x"9b",  x"22",  x"61",  x"f1",  x"3e",  x"01", -- 1098
         x"32",  x"eb",  x"f0",  x"32",  x"0e",  x"f1",  x"21",  x"bc", -- 10A0
         x"34",  x"22",  x"17",  x"f1",  x"21",  x"0b",  x"16",  x"22", -- 10A8
         x"15",  x"f1",  x"c9",  x"3a",  x"5f",  x"f1",  x"fe",  x"8b", -- 10B0
         x"ca",  x"bc",  x"30",  x"d8",  x"3a",  x"6f",  x"f1",  x"fe", -- 10B8
         x"18",  x"da",  x"e4",  x"2f",  x"fe",  x"2d",  x"d8",  x"fe", -- 10C0
         x"48",  x"da",  x"e4",  x"2f",  x"fe",  x"5d",  x"da",  x"01", -- 10C8
         x"31",  x"fe",  x"78",  x"da",  x"e4",  x"2f",  x"fe",  x"8d", -- 10D0
         x"da",  x"23",  x"31",  x"fe",  x"a0",  x"da",  x"f8",  x"30", -- 10D8
         x"3a",  x"eb",  x"f0",  x"fe",  x"04",  x"c8",  x"3e",  x"04", -- 10E0
         x"32",  x"eb",  x"f0",  x"21",  x"ae",  x"34",  x"22",  x"03", -- 10E8
         x"f1",  x"21",  x"07",  x"16",  x"22",  x"15",  x"f1",  x"c9", -- 10F0
         x"3a",  x"5f",  x"f1",  x"fe",  x"90",  x"d8",  x"c3",  x"e4", -- 10F8
         x"2f",  x"3a",  x"eb",  x"f0",  x"fe",  x"02",  x"c8",  x"32", -- 1100
         x"0f",  x"f1",  x"3a",  x"63",  x"f1",  x"fe",  x"ab",  x"c2", -- 1108
         x"e4",  x"2f",  x"21",  x"bc",  x"34",  x"22",  x"08",  x"f1", -- 1110
         x"21",  x"ae",  x"34",  x"22",  x"17",  x"f1",  x"3e",  x"02", -- 1118
         x"c3",  x"42",  x"31",  x"3a",  x"eb",  x"f0",  x"fe",  x"03", -- 1120
         x"c8",  x"32",  x"10",  x"f1",  x"3a",  x"66",  x"f1",  x"fe", -- 1128
         x"ab",  x"c2",  x"e4",  x"2f",  x"21",  x"bc",  x"34",  x"22", -- 1130
         x"03",  x"f1",  x"21",  x"ae",  x"34",  x"22",  x"08",  x"f1", -- 1138
         x"3e",  x"03",  x"32",  x"eb",  x"f0",  x"c9",  x"3e",  x"39", -- 1140
         x"32",  x"0b",  x"f1",  x"32",  x"ec",  x"f0",  x"cd",  x"36", -- 1148
         x"21",  x"3e",  x"ff",  x"32",  x"9d",  x"f1",  x"cd",  x"85", -- 1150
         x"21",  x"36",  x"a8",  x"23",  x"36",  x"b8",  x"23",  x"36", -- 1158
         x"b0",  x"21",  x"60",  x"70",  x"22",  x"77",  x"f1",  x"21", -- 1160
         x"b8",  x"b8",  x"22",  x"79",  x"f1",  x"21",  x"92",  x"92", -- 1168
         x"22",  x"5b",  x"f1",  x"21",  x"a2",  x"a2",  x"22",  x"5d", -- 1170
         x"f1",  x"21",  x"a5",  x"a5",  x"22",  x"67",  x"f1",  x"21", -- 1178
         x"9b",  x"9b",  x"22",  x"5f",  x"f1",  x"21",  x"ab",  x"ab", -- 1180
         x"22",  x"61",  x"f1",  x"22",  x"63",  x"f1",  x"22",  x"65", -- 1188
         x"f1",  x"21",  x"50",  x"60",  x"22",  x"69",  x"f1",  x"cd", -- 1190
         x"a5",  x"21",  x"21",  x"65",  x"75",  x"22",  x"87",  x"f1", -- 1198
         x"16",  x"46",  x"cd",  x"66",  x"1a",  x"11",  x"7b",  x"f1", -- 11A0
         x"cd",  x"82",  x"1a",  x"16",  x"3e",  x"cd",  x"66",  x"1a", -- 11A8
         x"11",  x"7f",  x"f1",  x"cd",  x"82",  x"1a",  x"21",  x"5d", -- 11B0
         x"5e",  x"22",  x"89",  x"f1",  x"21",  x"98",  x"34",  x"22", -- 11B8
         x"08",  x"f1",  x"af",  x"32",  x"eb",  x"f0",  x"3e",  x"01", -- 11C0
         x"32",  x"0f",  x"f1",  x"21",  x"e0",  x"17",  x"7e",  x"32", -- 11C8
         x"ef",  x"f0",  x"22",  x"06",  x"f1",  x"cd",  x"4a",  x"23", -- 11D0
         x"c3",  x"d9",  x"39",  x"cd",  x"f8",  x"31",  x"3a",  x"14", -- 11D8
         x"f1",  x"b7",  x"ca",  x"4c",  x"39",  x"3a",  x"6c",  x"f1", -- 11E0
         x"fe",  x"30",  x"da",  x"be",  x"37",  x"fe",  x"a0",  x"da", -- 11E8
         x"b6",  x"37",  x"cd",  x"d1",  x"32",  x"c3",  x"4c",  x"39", -- 11F0
         x"3a",  x"0f",  x"f1",  x"3d",  x"32",  x"0f",  x"f1",  x"c0", -- 11F8
         x"2a",  x"08",  x"f1",  x"7e",  x"fe",  x"2f",  x"c2",  x"84", -- 1200
         x"32",  x"3a",  x"a6",  x"f1",  x"fe",  x"58",  x"c2",  x"23", -- 1208
         x"32",  x"21",  x"94",  x"34",  x"22",  x"08",  x"f1",  x"3a", -- 1210
         x"ef",  x"f0",  x"3d",  x"32",  x"ef",  x"f0",  x"c2",  x"84", -- 1218
         x"32",  x"c1",  x"c9",  x"3a",  x"eb",  x"f0",  x"b7",  x"ca", -- 1220
         x"30",  x"32",  x"21",  x"82",  x"34",  x"c3",  x"84",  x"32", -- 1228
         x"23",  x"22",  x"08",  x"f1",  x"3a",  x"ef",  x"f0",  x"3d", -- 1230
         x"32",  x"ef",  x"f0",  x"11",  x"f3",  x"ff",  x"19",  x"c2", -- 1238
         x"84",  x"32",  x"2a",  x"06",  x"f1",  x"3a",  x"81",  x"f1", -- 1240
         x"fe",  x"58",  x"3e",  x"00",  x"c2",  x"51",  x"32",  x"3e", -- 1248
         x"10",  x"86",  x"32",  x"ef",  x"f0",  x"23",  x"7e",  x"fe", -- 1250
         x"ff",  x"c2",  x"5f",  x"32",  x"21",  x"e0",  x"17",  x"22", -- 1258
         x"06",  x"f1",  x"2a",  x"08",  x"f1",  x"7e",  x"fe",  x"2e", -- 1260
         x"ca",  x"76",  x"32",  x"3a",  x"5f",  x"f1",  x"c6",  x"08", -- 1268
         x"32",  x"5f",  x"f1",  x"c3",  x"84",  x"32",  x"3a",  x"5f", -- 1270
         x"f1",  x"c6",  x"f0",  x"32",  x"5f",  x"f1",  x"32",  x"60", -- 1278
         x"f1",  x"21",  x"94",  x"34",  x"23",  x"3a",  x"5f",  x"f1", -- 1280
         x"86",  x"32",  x"5f",  x"f1",  x"32",  x"60",  x"f1",  x"3a", -- 1288
         x"eb",  x"f0",  x"b7",  x"ca",  x"9d",  x"32",  x"7e",  x"11", -- 1290
         x"5b",  x"f1",  x"cd",  x"60",  x"1b",  x"23",  x"7e",  x"32", -- 1298
         x"0f",  x"f1",  x"23",  x"11",  x"7f",  x"f1",  x"cd",  x"4d", -- 12A0
         x"1b",  x"22",  x"08",  x"f1",  x"7e",  x"fe",  x"cc",  x"c0", -- 12A8
         x"23",  x"22",  x"08",  x"f1",  x"21",  x"82",  x"f1",  x"7e", -- 12B0
         x"b7",  x"ca",  x"c0",  x"32",  x"23",  x"c3",  x"b7",  x"32", -- 12B8
         x"3e",  x"08",  x"77",  x"11",  x"ef",  x"ff",  x"19",  x"7e", -- 12C0
         x"23",  x"77",  x"19",  x"7e",  x"c6",  x"f0",  x"23",  x"77", -- 12C8
         x"c9",  x"3a",  x"eb",  x"f0",  x"b7",  x"ca",  x"03",  x"33", -- 12D0
         x"3a",  x"a6",  x"f1",  x"fe",  x"58",  x"c8",  x"3a",  x"5b", -- 12D8
         x"f1",  x"fe",  x"50",  x"d0",  x"3a",  x"a6",  x"f1",  x"fe", -- 12E0
         x"58",  x"c8",  x"3e",  x"58",  x"32",  x"a6",  x"f1",  x"cd", -- 12E8
         x"e3",  x"0f",  x"21",  x"94",  x"34",  x"22",  x"08",  x"f1", -- 12F0
         x"3e",  x"30",  x"32",  x"ef",  x"f0",  x"3e",  x"01",  x"32", -- 12F8
         x"0f",  x"f1",  x"c9",  x"3a",  x"a6",  x"f1",  x"fe",  x"57", -- 1300
         x"c8",  x"fe",  x"4a",  x"c0",  x"3a",  x"fa",  x"f0",  x"fe", -- 1308
         x"49",  x"ca",  x"1d",  x"33",  x"3a",  x"5b",  x"f1",  x"fe", -- 1310
         x"8c",  x"d8",  x"c3",  x"7a",  x"33",  x"3a",  x"6b",  x"f1", -- 1318
         x"fe",  x"98",  x"da",  x"7a",  x"33",  x"fe",  x"a8",  x"d2", -- 1320
         x"7a",  x"33",  x"3a",  x"81",  x"f1",  x"b7",  x"ca",  x"3a", -- 1328
         x"33",  x"3a",  x"5b",  x"f1",  x"fe",  x"8c",  x"d8",  x"c3", -- 1330
         x"7a",  x"33",  x"3a",  x"5b",  x"f1",  x"47",  x"3a",  x"61", -- 1338
         x"f1",  x"90",  x"fe",  x"1f",  x"c0",  x"21",  x"8b",  x"8b", -- 1340
         x"22",  x"5b",  x"f1",  x"21",  x"9b",  x"9b",  x"22",  x"5d", -- 1348
         x"f1",  x"3e",  x"01",  x"32",  x"eb",  x"f0",  x"21",  x"00", -- 1350
         x"00",  x"22",  x"87",  x"f1",  x"21",  x"76",  x"34",  x"22", -- 1358
         x"08",  x"f1",  x"21",  x"0b",  x"16",  x"22",  x"15",  x"f1", -- 1360
         x"3e",  x"01",  x"32",  x"0f",  x"f1",  x"3e",  x"52",  x"32", -- 1368
         x"a6",  x"f1",  x"af",  x"32",  x"19",  x"f1",  x"cd",  x"e3", -- 1370
         x"0f",  x"c9",  x"af",  x"32",  x"19",  x"f1",  x"3e",  x"09", -- 1378
         x"32",  x"f5",  x"f0",  x"21",  x"a8",  x"a8",  x"22",  x"5b", -- 1380
         x"f1",  x"22",  x"5d",  x"f1",  x"3e",  x"57",  x"32",  x"a6", -- 1388
         x"f1",  x"af",  x"32",  x"14",  x"f1",  x"32",  x"eb",  x"f0", -- 1390
         x"cd",  x"e3",  x"0f",  x"21",  x"9a",  x"15",  x"11",  x"7b", -- 1398
         x"f1",  x"cd",  x"4d",  x"1b",  x"3a",  x"f9",  x"f0",  x"32", -- 13A0
         x"fa",  x"f0",  x"22",  x"15",  x"f1",  x"c9",  x"3e",  x"3a", -- 13A8
         x"cd",  x"75",  x"35",  x"21",  x"a3",  x"5d",  x"22",  x"83", -- 13B0
         x"f1",  x"21",  x"b3",  x"5e",  x"22",  x"85",  x"f1",  x"21", -- 13B8
         x"00",  x"00",  x"22",  x"7b",  x"f1",  x"3e",  x"09",  x"32", -- 13C0
         x"93",  x"f1",  x"32",  x"95",  x"f1",  x"21",  x"88",  x"98", -- 13C8
         x"22",  x"73",  x"f1",  x"22",  x"75",  x"f1",  x"21",  x"80", -- 13D0
         x"80",  x"22",  x"63",  x"f1",  x"21",  x"90",  x"90",  x"22", -- 13D8
         x"65",  x"f1",  x"cd",  x"41",  x"22",  x"cd",  x"57",  x"36", -- 13E0
         x"cd",  x"41",  x"22",  x"21",  x"17",  x"f1",  x"36",  x"33", -- 13E8
         x"11",  x"7f",  x"f1",  x"cd",  x"4d",  x"1b",  x"cd",  x"41", -- 13F0
         x"22",  x"21",  x"17",  x"f1",  x"36",  x"08",  x"cd",  x"88", -- 13F8
         x"36",  x"cd",  x"41",  x"22",  x"3a",  x"5f",  x"f1",  x"c6", -- 1400
         x"08",  x"32",  x"62",  x"f1",  x"3e",  x"01",  x"32",  x"13", -- 1408
         x"f1",  x"32",  x"0e",  x"f1",  x"af",  x"32",  x"14",  x"f1", -- 1410
         x"21",  x"00",  x"00",  x"22",  x"7f",  x"f1",  x"22",  x"81", -- 1418
         x"f1",  x"21",  x"ae",  x"16",  x"22",  x"a7",  x"f1",  x"cd", -- 1420
         x"98",  x"23",  x"3e",  x"05",  x"32",  x"93",  x"f1",  x"32", -- 1428
         x"95",  x"f1",  x"21",  x"6e",  x"5d",  x"22",  x"83",  x"f1", -- 1430
         x"21",  x"6f",  x"7a",  x"22",  x"85",  x"f1",  x"c3",  x"4c", -- 1438
         x"39",  x"3a",  x"82",  x"f1",  x"b7",  x"c2",  x"4c",  x"39", -- 1440
         x"3a",  x"88",  x"f1",  x"b7",  x"c8",  x"3a",  x"67",  x"f1", -- 1448
         x"c6",  x"08",  x"32",  x"62",  x"f1",  x"3a",  x"77",  x"f1", -- 1450
         x"c6",  x"08",  x"32",  x"72",  x"f1",  x"af",  x"32",  x"14", -- 1458
         x"f1",  x"21",  x"00",  x"00",  x"22",  x"87",  x"f1",  x"22", -- 1460
         x"89",  x"f1",  x"21",  x"ae",  x"16",  x"22",  x"a7",  x"f1", -- 1468
         x"cd",  x"98",  x"23",  x"c3",  x"4c",  x"39",  x"00",  x"00", -- 1470
         x"05",  x"64",  x"00",  x"fc",  x"05",  x"62",  x"00",  x"fc", -- 1478
         x"05",  x"63",  x"00",  x"fc",  x"05",  x"3e",  x"00",  x"fc", -- 1480
         x"05",  x"3f",  x"00",  x"fc",  x"05",  x"3e",  x"cc",  x"00", -- 1488
         x"fc",  x"05",  x"40",  x"2f",  x"00",  x"00",  x"01",  x"3e", -- 1490
         x"00",  x"00",  x"01",  x"3f",  x"00",  x"00",  x"01",  x"40", -- 1498
         x"2f",  x"00",  x"00",  x"01",  x"61",  x"00",  x"00",  x"01", -- 14A0
         x"62",  x"00",  x"00",  x"01",  x"63",  x"2f",  x"00",  x"00", -- 14A8
         x"01",  x"64",  x"00",  x"00",  x"01",  x"65",  x"00",  x"00", -- 14B0
         x"01",  x"66",  x"2f",  x"2e",  x"00",  x"00",  x"01",  x"64", -- 14B8
         x"00",  x"00",  x"01",  x"65",  x"00",  x"00",  x"01",  x"66", -- 14C0
         x"2f",  x"3e",  x"30",  x"cd",  x"75",  x"35",  x"cd",  x"41", -- 14C8
         x"22",  x"cd",  x"83",  x"36",  x"21",  x"4a",  x"5f",  x"22", -- 14D0
         x"83",  x"f1",  x"22",  x"0c",  x"f0",  x"21",  x"00",  x"00", -- 14D8
         x"22",  x"85",  x"f1",  x"22",  x"10",  x"f0",  x"cd",  x"05", -- 14E0
         x"36",  x"cd",  x"57",  x"36",  x"cd",  x"6d",  x"36",  x"cd", -- 14E8
         x"41",  x"22",  x"cd",  x"83",  x"36",  x"cd",  x"98",  x"36", -- 14F0
         x"c9",  x"3e",  x"30",  x"cd",  x"75",  x"35",  x"21",  x"4a", -- 14F8
         x"5f",  x"22",  x"83",  x"f1",  x"3a",  x"6b",  x"f1",  x"d6", -- 1500
         x"04",  x"32",  x"73",  x"f1",  x"c6",  x"0f",  x"32",  x"74", -- 1508
         x"f1",  x"3a",  x"5c",  x"f1",  x"32",  x"63",  x"f1",  x"32", -- 1510
         x"64",  x"f1",  x"cd",  x"c9",  x"36",  x"21",  x"3c",  x"4c", -- 1518
         x"22",  x"83",  x"f1",  x"22",  x"0c",  x"f0",  x"21",  x"4d", -- 1520
         x"85",  x"cd",  x"f8",  x"36",  x"c9",  x"3e",  x"30",  x"cd", -- 1528
         x"75",  x"35",  x"21",  x"3c",  x"4c",  x"22",  x"83",  x"f1", -- 1530
         x"21",  x"4d",  x"85",  x"22",  x"85",  x"f1",  x"3a",  x"6b", -- 1538
         x"f1",  x"d6",  x"03",  x"32",  x"74",  x"f1",  x"32",  x"76", -- 1540
         x"f1",  x"d6",  x"0f",  x"32",  x"73",  x"f1",  x"32",  x"75", -- 1548
         x"f1",  x"3a",  x"5b",  x"f1",  x"c6",  x"07",  x"21",  x"63", -- 1550
         x"f1",  x"77",  x"23",  x"77",  x"23",  x"c6",  x"0f",  x"77", -- 1558
         x"23",  x"77",  x"cd",  x"c9",  x"36",  x"21",  x"5d",  x"00", -- 1560
         x"22",  x"83",  x"f1",  x"22",  x"0c",  x"f0",  x"21",  x"5e", -- 1568
         x"00",  x"cd",  x"f8",  x"36",  x"c9",  x"32",  x"0b",  x"f1", -- 1570
         x"3a",  x"f2",  x"f0",  x"b7",  x"ca",  x"87",  x"35",  x"3e", -- 1578
         x"31",  x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"3e", -- 1580
         x"01",  x"32",  x"ec",  x"f0",  x"cd",  x"20",  x"21",  x"af", -- 1588
         x"32",  x"a4",  x"f1",  x"21",  x"70",  x"70",  x"22",  x"67", -- 1590
         x"f1",  x"21",  x"80",  x"80",  x"22",  x"5b",  x"f1",  x"22", -- 1598
         x"69",  x"f1",  x"22",  x"5f",  x"f1",  x"21",  x"90",  x"90", -- 15A0
         x"22",  x"5c",  x"f1",  x"22",  x"5d",  x"f1",  x"22",  x"61", -- 15A8
         x"f1",  x"21",  x"78",  x"78",  x"22",  x"63",  x"f1",  x"21", -- 15B0
         x"a0",  x"a0",  x"22",  x"6b",  x"f1",  x"21",  x"a8",  x"b8", -- 15B8
         x"22",  x"6d",  x"f1",  x"21",  x"50",  x"60",  x"22",  x"77", -- 15C0
         x"f1",  x"22",  x"79",  x"f1",  x"21",  x"78",  x"88",  x"22", -- 15C8
         x"73",  x"f1",  x"21",  x"20",  x"30",  x"22",  x"6f",  x"f1", -- 15D0
         x"22",  x"71",  x"f1",  x"21",  x"a3",  x"b3",  x"22",  x"7b", -- 15D8
         x"f1",  x"21",  x"6b",  x"6a",  x"22",  x"7d",  x"f1",  x"21", -- 15E0
         x"17",  x"f1",  x"36",  x"08",  x"11",  x"87",  x"f1",  x"cd", -- 15E8
         x"4d",  x"1b",  x"21",  x"70",  x"17",  x"11",  x"7f",  x"f1", -- 15F0
         x"cd",  x"4d",  x"1b",  x"21",  x"09",  x"09",  x"22",  x"8b", -- 15F8
         x"f1",  x"22",  x"8d",  x"f1",  x"c9",  x"0e",  x"08",  x"11", -- 1600
         x"09",  x"0c",  x"d5",  x"cd",  x"9f",  x"1a",  x"d1",  x"15", -- 1608
         x"c2",  x"2d",  x"36",  x"3a",  x"7d",  x"f1",  x"fe",  x"6d", -- 1610
         x"c2",  x"23",  x"36",  x"16",  x"0c",  x"21",  x"6b",  x"6a", -- 1618
         x"c3",  x"26",  x"36",  x"21",  x"6d",  x"6c",  x"22",  x"7d", -- 1620
         x"f1",  x"16",  x"08",  x"0d",  x"c8",  x"1d",  x"c2",  x"0a", -- 1628
         x"36",  x"3a",  x"83",  x"f1",  x"b7",  x"c2",  x"49",  x"36", -- 1630
         x"cd",  x"0b",  x"f0",  x"22",  x"83",  x"f1",  x"cd",  x"0f", -- 1638
         x"f0",  x"22",  x"85",  x"f1",  x"1e",  x"09",  x"c3",  x"0a", -- 1640
         x"36",  x"21",  x"00",  x"00",  x"22",  x"83",  x"f1",  x"22", -- 1648
         x"85",  x"f1",  x"1e",  x"03",  x"c3",  x"0a",  x"36",  x"21", -- 1650
         x"80",  x"f3",  x"22",  x"87",  x"f1",  x"21",  x"82",  x"81", -- 1658
         x"22",  x"89",  x"f1",  x"21",  x"09",  x"09",  x"22",  x"97", -- 1660
         x"f1",  x"22",  x"99",  x"f1",  x"c9",  x"21",  x"6a",  x"6b", -- 1668
         x"22",  x"7d",  x"f1",  x"21",  x"05",  x"05",  x"22",  x"8b", -- 1670
         x"f1",  x"22",  x"8d",  x"f1",  x"21",  x"a8",  x"a8",  x"22", -- 1678
         x"6b",  x"f1",  x"c9",  x"21",  x"17",  x"f1",  x"36",  x"09", -- 1680
         x"11",  x"87",  x"f1",  x"cd",  x"4d",  x"1b",  x"21",  x"05", -- 1688
         x"05",  x"22",  x"97",  x"f1",  x"22",  x"99",  x"f1",  x"c9", -- 1690
         x"3a",  x"f2",  x"f0",  x"b7",  x"c0",  x"21",  x"a0",  x"b0", -- 1698
         x"22",  x"6b",  x"f1",  x"22",  x"6d",  x"f1",  x"3e",  x"80", -- 16A0
         x"32",  x"5c",  x"f1",  x"cd",  x"a5",  x"21",  x"cd",  x"41", -- 16A8
         x"22",  x"c3",  x"16",  x"3c",  x"3a",  x"6b",  x"f1",  x"fe", -- 16B0
         x"c8",  x"d2",  x"c2",  x"36",  x"cd",  x"9f",  x"1a",  x"c3", -- 16B8
         x"64",  x"39",  x"cd",  x"20",  x"21",  x"cd",  x"9f",  x"1a", -- 16C0
         x"c9",  x"cd",  x"41",  x"22",  x"cd",  x"57",  x"36",  x"cd", -- 16C8
         x"41",  x"22",  x"21",  x"17",  x"f1",  x"36",  x"33",  x"11", -- 16D0
         x"7f",  x"f1",  x"cd",  x"4d",  x"1b",  x"cd",  x"41",  x"22", -- 16D8
         x"21",  x"70",  x"17",  x"11",  x"7f",  x"f1",  x"cd",  x"4d", -- 16E0
         x"1b",  x"21",  x"17",  x"f1",  x"36",  x"08",  x"cd",  x"88", -- 16E8
         x"36",  x"cd",  x"41",  x"22",  x"cd",  x"83",  x"36",  x"c9", -- 16F0
         x"22",  x"85",  x"f1",  x"22",  x"10",  x"f0",  x"21",  x"78", -- 16F8
         x"88",  x"22",  x"73",  x"f1",  x"22",  x"75",  x"f1",  x"21", -- 1700
         x"70",  x"70",  x"22",  x"63",  x"f1",  x"21",  x"80",  x"80", -- 1708
         x"22",  x"65",  x"f1",  x"cd",  x"05",  x"36",  x"cd",  x"6d", -- 1710
         x"36",  x"cd",  x"41",  x"22",  x"cd",  x"98",  x"36",  x"c9", -- 1718
         x"cd",  x"31",  x"3f",  x"3e",  x"31",  x"32",  x"0b",  x"f1", -- 1720
         x"cd",  x"36",  x"21",  x"cd",  x"2c",  x"22",  x"cd",  x"13", -- 1728
         x"22",  x"3e",  x"01",  x"32",  x"1a",  x"f1",  x"cd",  x"85", -- 1730
         x"21",  x"36",  x"70",  x"cd",  x"95",  x"21",  x"3e",  x"a8", -- 1738
         x"02",  x"cd",  x"a5",  x"21",  x"36",  x"93",  x"c3",  x"4c", -- 1740
         x"39",  x"3e",  x"32",  x"32",  x"0b",  x"f1",  x"32",  x"ec", -- 1748
         x"f0",  x"3e",  x"93",  x"32",  x"ff",  x"f0",  x"cd",  x"d6", -- 1750
         x"21",  x"cd",  x"2c",  x"22",  x"cd",  x"80",  x"22",  x"c3", -- 1758
         x"4c",  x"39",  x"21",  x"80",  x"f1",  x"22",  x"08",  x"f0", -- 1760
         x"01",  x"50",  x"06",  x"cd",  x"20",  x"22",  x"c3",  x"a6", -- 1768
         x"3e",  x"3e",  x"33",  x"32",  x"0b",  x"f1",  x"32",  x"ec", -- 1770
         x"f0",  x"cd",  x"36",  x"21",  x"3e",  x"ff",  x"32",  x"9d", -- 1778
         x"f1",  x"cd",  x"85",  x"21",  x"21",  x"90",  x"a0",  x"22", -- 1780
         x"77",  x"f1",  x"cd",  x"95",  x"21",  x"21",  x"a8",  x"a8", -- 1788
         x"22",  x"67",  x"f1",  x"cd",  x"a5",  x"21",  x"21",  x"65", -- 1790
         x"75",  x"22",  x"87",  x"f1",  x"cd",  x"4a",  x"23",  x"c3", -- 1798
         x"ad",  x"39",  x"3a",  x"14",  x"f1",  x"b7",  x"ca",  x"4c", -- 17A0
         x"39",  x"3a",  x"6c",  x"f1",  x"fe",  x"50",  x"da",  x"be", -- 17A8
         x"37",  x"fe",  x"d8",  x"d2",  x"be",  x"37",  x"3e",  x"01", -- 17B0
         x"32",  x"9c",  x"f1",  x"c3",  x"c7",  x"37",  x"af",  x"32", -- 17B8
         x"9c",  x"f1",  x"3e",  x"01",  x"32",  x"9b",  x"f1",  x"3a", -- 17C0
         x"a6",  x"f1",  x"fe",  x"4a",  x"c2",  x"de",  x"37",  x"3a", -- 17C8
         x"9b",  x"f1",  x"b7",  x"ca",  x"e8",  x"37",  x"3a",  x"fa", -- 17D0
         x"f0",  x"fe",  x"46",  x"c2",  x"e5",  x"37",  x"3a",  x"9c", -- 17D8
         x"f1",  x"b7",  x"c2",  x"f0",  x"37",  x"c3",  x"a6",  x"3e", -- 17E0
         x"3e",  x"01",  x"32",  x"9b",  x"f1",  x"c3",  x"a6",  x"3e", -- 17E8
         x"2a",  x"6b",  x"f1",  x"3a",  x"77",  x"f1",  x"c6",  x"08", -- 17F0
         x"bc",  x"d2",  x"19",  x"38",  x"c6",  x"10",  x"bc",  x"da", -- 17F8
         x"19",  x"38",  x"af",  x"32",  x"19",  x"f1",  x"32",  x"9b", -- 1800
         x"f1",  x"3e",  x"01",  x"32",  x"13",  x"f1",  x"3e",  x"53", -- 1808
         x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"c3",  x"a6", -- 1810
         x"3e",  x"3a",  x"6b",  x"f1",  x"fe",  x"a0",  x"d2",  x"49", -- 1818
         x"38",  x"01",  x"0f",  x"04",  x"21",  x"6b",  x"f1",  x"79", -- 1820
         x"86",  x"77",  x"23",  x"05",  x"c2",  x"27",  x"38",  x"3e", -- 1828
         x"01",  x"32",  x"f5",  x"f0",  x"21",  x"9b",  x"15",  x"22", -- 1830
         x"15",  x"f1",  x"af",  x"32",  x"14",  x"f1",  x"3e",  x"57", -- 1838
         x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"c3",  x"4c", -- 1840
         x"39",  x"01",  x"f1",  x"04",  x"c3",  x"24",  x"38",  x"3e", -- 1848
         x"34",  x"32",  x"0b",  x"f1",  x"32",  x"ec",  x"f0",  x"cd", -- 1850
         x"36",  x"21",  x"cd",  x"85",  x"21",  x"36",  x"60",  x"23", -- 1858
         x"36",  x"d0",  x"23",  x"36",  x"28",  x"23",  x"36",  x"90", -- 1860
         x"cd",  x"95",  x"21",  x"11",  x"9e",  x"f1",  x"3e",  x"20", -- 1868
         x"02",  x"12",  x"03",  x"13",  x"3e",  x"1e",  x"02",  x"12", -- 1870
         x"03",  x"13",  x"3e",  x"30",  x"02",  x"12",  x"03",  x"13", -- 1878
         x"3e",  x"25",  x"02",  x"12",  x"cd",  x"a5",  x"21",  x"06", -- 1880
         x"04",  x"36",  x"46",  x"23",  x"05",  x"c2",  x"89",  x"38", -- 1888
         x"cd",  x"9f",  x"1a",  x"cd",  x"75",  x"23",  x"c3",  x"96", -- 1890
         x"39",  x"3e",  x"36",  x"32",  x"0b",  x"f1",  x"32",  x"ec", -- 1898
         x"f0",  x"cd",  x"36",  x"21",  x"cd",  x"85",  x"21",  x"cd", -- 18A0
         x"95",  x"21",  x"cd",  x"a5",  x"21",  x"21",  x"82",  x"f1", -- 18A8
         x"cd",  x"4c",  x"22",  x"c3",  x"4c",  x"39",  x"3e",  x"37", -- 18B0
         x"32",  x"0b",  x"f1",  x"32",  x"ec",  x"f0",  x"3e",  x"54", -- 18B8
         x"32",  x"ff",  x"f0",  x"cd",  x"d6",  x"21",  x"cd",  x"af", -- 18C0
         x"22",  x"cd",  x"80",  x"22",  x"23",  x"cd",  x"4c",  x"22", -- 18C8
         x"c3",  x"4c",  x"39",  x"3e",  x"35",  x"32",  x"0b",  x"f1", -- 18D0
         x"32",  x"ec",  x"f0",  x"cd",  x"36",  x"21",  x"cd",  x"85", -- 18D8
         x"21",  x"21",  x"d2",  x"e2",  x"22",  x"6f",  x"f1",  x"3e", -- 18E0
         x"c0",  x"32",  x"72",  x"f1",  x"21",  x"d0",  x"e4",  x"22", -- 18E8
         x"73",  x"f1",  x"21",  x"d7",  x"e7",  x"22",  x"75",  x"f1", -- 18F0
         x"22",  x"77",  x"f1",  x"cd",  x"95",  x"21",  x"3e",  x"9d", -- 18F8
         x"02",  x"03",  x"02",  x"03",  x"03",  x"3e",  x"a2",  x"02", -- 1900
         x"03",  x"3e",  x"a8",  x"02",  x"03",  x"02",  x"03",  x"3e", -- 1908
         x"89",  x"02",  x"03",  x"02",  x"03",  x"3e",  x"99",  x"02", -- 1910
         x"03",  x"02",  x"cd",  x"a5",  x"21",  x"21",  x"43",  x"63", -- 1918
         x"22",  x"7f",  x"f1",  x"3e",  x"0a",  x"32",  x"82",  x"f1", -- 1920
         x"21",  x"84",  x"84",  x"22",  x"83",  x"f1",  x"21",  x"3c", -- 1928
         x"4c",  x"22",  x"85",  x"f1",  x"21",  x"4d",  x"85",  x"22", -- 1930
         x"87",  x"f1",  x"cd",  x"9f",  x"1a",  x"21",  x"f2",  x"16", -- 1938
         x"22",  x"a7",  x"f1",  x"21",  x"3d",  x"17",  x"22",  x"08", -- 1940
         x"f1",  x"c3",  x"4c",  x"39",  x"3a",  x"13",  x"f1",  x"b7", -- 1948
         x"c2",  x"6e",  x"39",  x"3a",  x"f8",  x"f0",  x"b7",  x"ca", -- 1950
         x"64",  x"39",  x"3d",  x"32",  x"f8",  x"f0",  x"c2",  x"64", -- 1958
         x"39",  x"32",  x"8a",  x"f1",  x"3a",  x"f5",  x"f0",  x"3d", -- 1960
         x"32",  x"f5",  x"f0",  x"ca",  x"5d",  x"3c",  x"3a",  x"a4", -- 1968
         x"f1",  x"b7",  x"c2",  x"e5",  x"21",  x"3a",  x"0b",  x"f1", -- 1970
         x"d6",  x"30",  x"87",  x"5f",  x"16",  x"00",  x"21",  x"38", -- 1978
         x"1a",  x"19",  x"5e",  x"23",  x"56",  x"eb",  x"22",  x"05", -- 1980
         x"f0",  x"cd",  x"03",  x"f0",  x"3a",  x"0e",  x"f1",  x"3d", -- 1988
         x"32",  x"0e",  x"f1",  x"cc",  x"75",  x"23",  x"3a",  x"0f", -- 1990
         x"f1",  x"3d",  x"32",  x"0f",  x"f1",  x"cc",  x"86",  x"23", -- 1998
         x"c3",  x"69",  x"3a",  x"3a",  x"0e",  x"f1",  x"3d",  x"32", -- 19A0
         x"0e",  x"f1",  x"cc",  x"4a",  x"23",  x"3a",  x"77",  x"f1", -- 19A8
         x"fe",  x"54",  x"ca",  x"ba",  x"39",  x"fe",  x"b4",  x"c2", -- 19B0
         x"69",  x"3a",  x"3a",  x"9d",  x"f1",  x"2f",  x"3c",  x"32", -- 19B8
         x"9d",  x"f1",  x"cd",  x"4f",  x"23",  x"c3",  x"ad",  x"39", -- 19C0
         x"3a",  x"eb",  x"f0",  x"b7",  x"c2",  x"69",  x"3a",  x"3a", -- 19C8
         x"0e",  x"f1",  x"3d",  x"32",  x"0e",  x"f1",  x"cc",  x"4a", -- 19D0
         x"23",  x"3a",  x"77",  x"f1",  x"fe",  x"2c",  x"ca",  x"e6", -- 19D8
         x"39",  x"fe",  x"84",  x"c2",  x"69",  x"3a",  x"3a",  x"9d", -- 19E0
         x"f1",  x"2f",  x"3c",  x"32",  x"9d",  x"f1",  x"cd",  x"4f", -- 19E8
         x"23",  x"c3",  x"d9",  x"39",  x"3a",  x"0e",  x"f1",  x"b7", -- 19F0
         x"c2",  x"25",  x"3a",  x"3a",  x"e7",  x"f0",  x"3d",  x"32", -- 19F8
         x"e7",  x"f0",  x"c2",  x"46",  x"3a",  x"2a",  x"06",  x"f1", -- 1A00
         x"23",  x"22",  x"06",  x"f1",  x"7e",  x"fe",  x"ff",  x"ca", -- 1A08
         x"1f",  x"3a",  x"c6",  x"01",  x"32",  x"e7",  x"f0",  x"3e", -- 1A10
         x"01",  x"32",  x"0e",  x"f1",  x"c3",  x"46",  x"3a",  x"21", -- 1A18
         x"e0",  x"17",  x"c3",  x"09",  x"3a",  x"3a",  x"63",  x"f1", -- 1A20
         x"c6",  x"04",  x"32",  x"63",  x"f1",  x"fe",  x"a7",  x"da", -- 1A28
         x"46",  x"3a",  x"af",  x"32",  x"0e",  x"f1",  x"3a",  x"72", -- 1A30
         x"f1",  x"c6",  x"08",  x"32",  x"73",  x"f1",  x"3a",  x"62", -- 1A38
         x"f1",  x"c6",  x"06",  x"32",  x"63",  x"f1",  x"3a",  x"0f", -- 1A40
         x"f1",  x"3d",  x"32",  x"0f",  x"f1",  x"cc",  x"98",  x"23", -- 1A48
         x"3a",  x"0b",  x"f1",  x"fe",  x"35",  x"c2",  x"69",  x"3a", -- 1A50
         x"3a",  x"a5",  x"f1",  x"b7",  x"ca",  x"69",  x"3a",  x"3a", -- 1A58
         x"f6",  x"f0",  x"3d",  x"32",  x"f6",  x"f0",  x"cc",  x"f8", -- 1A60
         x"22",  x"cd",  x"9f",  x"1a",  x"3a",  x"14",  x"f1",  x"b7", -- 1A68
         x"ca",  x"8c",  x"3a",  x"3a",  x"0b",  x"f1",  x"fe",  x"3b", -- 1A70
         x"ca",  x"8c",  x"3a",  x"3a",  x"6c",  x"f1",  x"fe",  x"f0", -- 1A78
         x"da",  x"8c",  x"3a",  x"3a",  x"0b",  x"f1",  x"fe",  x"37", -- 1A80
         x"cc",  x"b5",  x"21",  x"c9",  x"3a",  x"0b",  x"f1",  x"d6", -- 1A88
         x"31",  x"87",  x"5f",  x"16",  x"00",  x"21",  x"50",  x"1a", -- 1A90
         x"19",  x"5e",  x"23",  x"56",  x"eb",  x"22",  x"05",  x"f0", -- 1A98
         x"cd",  x"03",  x"f0",  x"11",  x"5f",  x"f1",  x"21",  x"9e", -- 1AA0
         x"f1",  x"06",  x"04",  x"1a",  x"fe",  x"a5",  x"da",  x"b3", -- 1AA8
         x"3a",  x"7e",  x"12",  x"23",  x"13",  x"05",  x"c2",  x"ab", -- 1AB0
         x"3a",  x"3a",  x"14",  x"f1",  x"b7",  x"ca",  x"e3",  x"3a", -- 1AB8
         x"06",  x"05",  x"21",  x"6f",  x"f1",  x"11",  x"5f",  x"f1", -- 1AC0
         x"05",  x"ca",  x"e3",  x"3a",  x"3a",  x"6b",  x"f1",  x"be", -- 1AC8
         x"d2",  x"e6",  x"3a",  x"c6",  x"10",  x"be",  x"da",  x"e6", -- 1AD0
         x"3a",  x"21",  x"5b",  x"f1",  x"1a",  x"c6",  x"0c",  x"be", -- 1AD8
         x"d2",  x"29",  x"3e",  x"c3",  x"a6",  x"3e",  x"23",  x"13", -- 1AE0
         x"c3",  x"c8",  x"3a",  x"3a",  x"0b",  x"f1",  x"fe",  x"36", -- 1AE8
         x"ca",  x"a6",  x"3e",  x"3a",  x"1a",  x"f1",  x"b7",  x"ca", -- 1AF0
         x"a6",  x"3e",  x"3a",  x"14",  x"f1",  x"b7",  x"ca",  x"a6", -- 1AF8
         x"3e",  x"21",  x"6c",  x"f1",  x"3a",  x"a3",  x"f1",  x"be", -- 1B00
         x"d2",  x"23",  x"3b",  x"af",  x"cd",  x"07",  x"f0",  x"3a", -- 1B08
         x"1a",  x"f1",  x"3d",  x"32",  x"1a",  x"f1",  x"fe",  x"02", -- 1B10
         x"ca",  x"62",  x"37",  x"fe",  x"01",  x"cc",  x"13",  x"22", -- 1B18
         x"c3",  x"a6",  x"3e",  x"3a",  x"a6",  x"f1",  x"fe",  x"4a", -- 1B20
         x"ca",  x"41",  x"3b",  x"fe",  x"47",  x"c2",  x"a6",  x"3e", -- 1B28
         x"3a",  x"a0",  x"f1",  x"be",  x"d2",  x"a6",  x"3e",  x"3a", -- 1B30
         x"a1",  x"f1",  x"be",  x"da",  x"a6",  x"3e",  x"c3",  x"2c", -- 1B38
         x"3e",  x"3a",  x"fa",  x"f0",  x"fe",  x"47",  x"c2",  x"64", -- 1B40
         x"3b",  x"3a",  x"9f",  x"f1",  x"be",  x"d2",  x"a6",  x"3e", -- 1B48
         x"3a",  x"a2",  x"f1",  x"be",  x"da",  x"a6",  x"3e",  x"af", -- 1B50
         x"32",  x"14",  x"f1",  x"21",  x"15",  x"16",  x"22",  x"15", -- 1B58
         x"f1",  x"c3",  x"a6",  x"3e",  x"fe",  x"49",  x"c2",  x"a6", -- 1B60
         x"3e",  x"3a",  x"9e",  x"f1",  x"be",  x"d2",  x"a6",  x"3e", -- 1B68
         x"c3",  x"37",  x"3b",  x"3a",  x"14",  x"f1",  x"b7",  x"ca", -- 1B70
         x"a6",  x"3e",  x"3a",  x"0e",  x"f1",  x"b7",  x"ca",  x"eb", -- 1B78
         x"3a",  x"21",  x"73",  x"f1",  x"3a",  x"6b",  x"f1",  x"be", -- 1B80
         x"d2",  x"eb",  x"3a",  x"c6",  x"10",  x"be",  x"da",  x"eb", -- 1B88
         x"3a",  x"21",  x"5b",  x"f1",  x"3a",  x"63",  x"f1",  x"c6", -- 1B90
         x"0c",  x"be",  x"da",  x"eb",  x"3a",  x"af",  x"32",  x"0e", -- 1B98
         x"f1",  x"3a",  x"72",  x"f1",  x"c6",  x"08",  x"32",  x"73", -- 1BA0
         x"f1",  x"3a",  x"62",  x"f1",  x"c6",  x"06",  x"32",  x"63", -- 1BA8
         x"f1",  x"c3",  x"2c",  x"3e",  x"3a",  x"14",  x"f1",  x"b7", -- 1BB0
         x"ca",  x"4c",  x"39",  x"3a",  x"9b",  x"f1",  x"b7",  x"c2", -- 1BB8
         x"e3",  x"3b",  x"3a",  x"a5",  x"f1",  x"b7",  x"c2",  x"4c", -- 1BC0
         x"39",  x"21",  x"6c",  x"f1",  x"3a",  x"74",  x"f1",  x"c6", -- 1BC8
         x"1a",  x"be",  x"d2",  x"4c",  x"39",  x"3e",  x"01",  x"32", -- 1BD0
         x"a5",  x"f1",  x"21",  x"5f",  x"17",  x"22",  x"08",  x"f1", -- 1BD8
         x"c3",  x"4c",  x"39",  x"21",  x"72",  x"f1",  x"3a",  x"6b", -- 1BE0
         x"f1",  x"c6",  x"16",  x"be",  x"da",  x"a6",  x"3e",  x"3a", -- 1BE8
         x"a6",  x"f1",  x"fe",  x"59",  x"ca",  x"fd",  x"3b",  x"cd", -- 1BF0
         x"c4",  x"22",  x"c3",  x"5d",  x"3c",  x"21",  x"ae",  x"16", -- 1BF8
         x"22",  x"a7",  x"f1",  x"af",  x"32",  x"9b",  x"f1",  x"32", -- 1C00
         x"a5",  x"f1",  x"21",  x"09",  x"09",  x"22",  x"93",  x"f1", -- 1C08
         x"cd",  x"98",  x"23",  x"c3",  x"69",  x"3a",  x"06",  x"04", -- 1C10
         x"11",  x"6b",  x"f1",  x"1a",  x"3c",  x"12",  x"13",  x"05", -- 1C18
         x"c2",  x"1b",  x"3c",  x"3e",  x"0b",  x"32",  x"f5",  x"f0", -- 1C20
         x"3e",  x"34",  x"32",  x"fa",  x"f0",  x"21",  x"af",  x"15", -- 1C28
         x"11",  x"7b",  x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"15", -- 1C30
         x"f1",  x"c3",  x"6e",  x"39",  x"3a",  x"a6",  x"f1",  x"fe", -- 1C38
         x"46",  x"c2",  x"4a",  x"3c",  x"21",  x"c4",  x"44",  x"c3", -- 1C40
         x"60",  x"3c",  x"3a",  x"a4",  x"f1",  x"b7",  x"ca",  x"57", -- 1C48
         x"3c",  x"21",  x"6d",  x"16",  x"c3",  x"60",  x"3c",  x"21", -- 1C50
         x"b0",  x"15",  x"c3",  x"60",  x"3c",  x"2a",  x"15",  x"f1", -- 1C58
         x"7e",  x"fe",  x"2e",  x"ca",  x"fa",  x"3c",  x"fe",  x"2f", -- 1C60
         x"ca",  x"3c",  x"3c",  x"01",  x"02",  x"04",  x"11",  x"6b", -- 1C68
         x"f1",  x"1a",  x"86",  x"12",  x"13",  x"05",  x"c2",  x"71", -- 1C70
         x"3c",  x"23",  x"0d",  x"ca",  x"86",  x"3c",  x"06",  x"04", -- 1C78
         x"11",  x"5b",  x"f1",  x"c3",  x"71",  x"3c",  x"7e",  x"32", -- 1C80
         x"f5",  x"f0",  x"23",  x"11",  x"7b",  x"f1",  x"cd",  x"4d", -- 1C88
         x"1b",  x"22",  x"15",  x"f1",  x"7e",  x"fe",  x"cc",  x"c2", -- 1C90
         x"bc",  x"3c",  x"23",  x"3a",  x"6b",  x"f1",  x"86",  x"32", -- 1C98
         x"7a",  x"f1",  x"23",  x"3a",  x"5d",  x"f1",  x"86",  x"32", -- 1CA0
         x"6a",  x"f1",  x"23",  x"7e",  x"32",  x"f8",  x"f0",  x"23", -- 1CA8
         x"11",  x"8a",  x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"15", -- 1CB0
         x"f1",  x"c3",  x"6e",  x"39",  x"3a",  x"f9",  x"f0",  x"32", -- 1CB8
         x"fa",  x"f0",  x"fe",  x"31",  x"ca",  x"e8",  x"3c",  x"fe", -- 1CC0
         x"01",  x"ca",  x"f4",  x"3c",  x"2b",  x"11",  x"24",  x"16", -- 1CC8
         x"7a",  x"bc",  x"c2",  x"6e",  x"39",  x"7b",  x"bd",  x"c2", -- 1CD0
         x"6e",  x"39",  x"3a",  x"6b",  x"f1",  x"d6",  x"0c",  x"32", -- 1CD8
         x"74",  x"f1",  x"cd",  x"10",  x"21",  x"c3",  x"6e",  x"39", -- 1CE0
         x"21",  x"09",  x"09",  x"22",  x"8b",  x"f1",  x"22",  x"8d", -- 1CE8
         x"f1",  x"c3",  x"6e",  x"39",  x"21",  x"05",  x"05",  x"c3", -- 1CF0
         x"eb",  x"3c",  x"3a",  x"a4",  x"f1",  x"b7",  x"c2",  x"f3", -- 1CF8
         x"21",  x"3e",  x"01",  x"32",  x"19",  x"f1",  x"32",  x"13", -- 1D00
         x"f1",  x"3a",  x"a6",  x"f1",  x"fe",  x"52",  x"ca",  x"34", -- 1D08
         x"3d",  x"fe",  x"4c",  x"ca",  x"1e",  x"3d",  x"3e",  x"53", -- 1D10
         x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"3a",  x"0b", -- 1D18
         x"f1",  x"fe",  x"35",  x"c2",  x"34",  x"3d",  x"3a",  x"9b", -- 1D20
         x"f1",  x"b7",  x"c2",  x"34",  x"3d",  x"af",  x"32",  x"13", -- 1D28
         x"f1",  x"c3",  x"16",  x"3c",  x"3a",  x"14",  x"f1",  x"b7", -- 1D30
         x"c2",  x"4c",  x"39",  x"cd",  x"2c",  x"24",  x"c3",  x"19", -- 1D38
         x"3f",  x"af",  x"32",  x"19",  x"f1",  x"3a",  x"9b",  x"f1", -- 1D40
         x"b7",  x"c2",  x"63",  x"3d",  x"3a",  x"9d",  x"f1",  x"fe", -- 1D48
         x"01",  x"c2",  x"63",  x"3d",  x"2f",  x"3c",  x"32",  x"9d", -- 1D50
         x"f1",  x"3a",  x"0f",  x"f1",  x"2f",  x"3c",  x"c6",  x"50", -- 1D58
         x"32",  x"0f",  x"f1",  x"3a",  x"fa",  x"f0",  x"fe",  x"46", -- 1D60
         x"ca",  x"8c",  x"3d",  x"fe",  x"34",  x"ca",  x"ac",  x"3d", -- 1D68
         x"fe",  x"35",  x"ca",  x"b2",  x"3d",  x"fe",  x"36",  x"ca", -- 1D70
         x"ac",  x"3d",  x"fe",  x"37",  x"ca",  x"b2",  x"3d",  x"fe", -- 1D78
         x"3b",  x"ca",  x"b2",  x"3d",  x"3e",  x"01",  x"32",  x"19", -- 1D80
         x"f1",  x"c3",  x"4c",  x"39",  x"3a",  x"a6",  x"f1",  x"fe", -- 1D88
         x"53",  x"ca",  x"fa",  x"3c",  x"fe",  x"42",  x"ca",  x"07", -- 1D90
         x"3e",  x"fe",  x"59",  x"ca",  x"fe",  x"3d",  x"21",  x"ef", -- 1D98
         x"15",  x"22",  x"15",  x"f1",  x"3e",  x"01",  x"32",  x"f5", -- 1DA0
         x"f0",  x"c3",  x"6e",  x"39",  x"3a",  x"fb",  x"f0",  x"c3", -- 1DA8
         x"bb",  x"3d",  x"3a",  x"fc",  x"f0",  x"c3",  x"bb",  x"3d", -- 1DB0
         x"3a",  x"fd",  x"f0",  x"06",  x"04",  x"4f",  x"11",  x"6b", -- 1DB8
         x"f1",  x"1a",  x"81",  x"12",  x"13",  x"05",  x"c2",  x"c1", -- 1DC0
         x"3d",  x"3e",  x"4a",  x"32",  x"fa",  x"f0",  x"21",  x"ea", -- 1DC8
         x"15",  x"11",  x"7b",  x"f1",  x"cd",  x"4d",  x"1b",  x"22", -- 1DD0
         x"15",  x"f1",  x"3e",  x"0b",  x"32",  x"f5",  x"f0",  x"3a", -- 1DD8
         x"a6",  x"f1",  x"fe",  x"53",  x"c2",  x"f0",  x"3d",  x"21", -- 1DE0
         x"67",  x"16",  x"22",  x"15",  x"f1",  x"c3",  x"6e",  x"39", -- 1DE8
         x"fe",  x"59",  x"c2",  x"6e",  x"39",  x"21",  x"c2",  x"15", -- 1DF0
         x"22",  x"15",  x"f1",  x"c3",  x"6e",  x"39",  x"21",  x"c6", -- 1DF8
         x"15",  x"22",  x"15",  x"f1",  x"c3",  x"5d",  x"3c",  x"21", -- 1E00
         x"e1",  x"15",  x"22",  x"15",  x"f1",  x"c3",  x"5d",  x"3c", -- 1E08
         x"3e",  x"0b",  x"32",  x"f5",  x"f0",  x"3e",  x"3b",  x"32", -- 1E10
         x"fa",  x"f0",  x"21",  x"81",  x"16",  x"11",  x"7b",  x"f1", -- 1E18
         x"cd",  x"4d",  x"1b",  x"22",  x"15",  x"f1",  x"c3",  x"4c", -- 1E20
         x"39",  x"3e",  x"20",  x"12",  x"af",  x"32",  x"19",  x"f1", -- 1E28
         x"32",  x"13",  x"f1",  x"32",  x"14",  x"f1",  x"3a",  x"a6", -- 1E30
         x"f1",  x"fe",  x"47",  x"ca",  x"98",  x"3e",  x"3a",  x"fa", -- 1E38
         x"f0",  x"fe",  x"4a",  x"ca",  x"98",  x"3e",  x"fe",  x"46", -- 1E40
         x"ca",  x"98",  x"3e",  x"fe",  x"49",  x"ca",  x"56",  x"3e", -- 1E48
         x"21",  x"1d",  x"16",  x"c3",  x"8a",  x"3e",  x"3a",  x"6b", -- 1E50
         x"f1",  x"c6",  x"1a",  x"32",  x"74",  x"f1",  x"11",  x"f9", -- 1E58
         x"26",  x"01",  x"02",  x"04",  x"21",  x"6b",  x"f1",  x"7a", -- 1E60
         x"86",  x"77",  x"23",  x"05",  x"c2",  x"67",  x"3e",  x"21", -- 1E68
         x"5b",  x"f1",  x"06",  x"04",  x"53",  x"0d",  x"c2",  x"67", -- 1E70
         x"3e",  x"3e",  x"01",  x"32",  x"f5",  x"f0",  x"cd",  x"10", -- 1E78
         x"21",  x"21",  x"24",  x"16",  x"11",  x"7b",  x"f1",  x"cd", -- 1E80
         x"4d",  x"1b",  x"22",  x"15",  x"f1",  x"3e",  x"4b",  x"32", -- 1E88
         x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"c3",  x"6e",  x"39", -- 1E90
         x"3a",  x"6b",  x"f1",  x"c6",  x"0f",  x"32",  x"74",  x"f1", -- 1E98
         x"11",  x"f5",  x"1b",  x"c3",  x"61",  x"3e",  x"cd",  x"b6", -- 1EA0
         x"20",  x"ca",  x"4c",  x"39",  x"4f",  x"3a",  x"14",  x"f1", -- 1EA8
         x"b7",  x"ca",  x"4c",  x"39",  x"3a",  x"a6",  x"f1",  x"fe", -- 1EB0
         x"52",  x"ca",  x"1e",  x"45",  x"3a",  x"19",  x"f1",  x"b7", -- 1EB8
         x"ca",  x"04",  x"3f",  x"79",  x"fe",  x"47",  x"c2",  x"cf", -- 1EC0
         x"3e",  x"cd",  x"10",  x"3f",  x"c3",  x"16",  x"3c",  x"fe", -- 1EC8
         x"4c",  x"c2",  x"da",  x"3e",  x"cd",  x"10",  x"3f",  x"c3", -- 1ED0
         x"10",  x"3e",  x"fe",  x"59",  x"c2",  x"e7",  x"3e",  x"3a", -- 1ED8
         x"0b",  x"f1",  x"fe",  x"39",  x"c2",  x"0a",  x"3f",  x"fe", -- 1EE0
         x"53",  x"ca",  x"0a",  x"3f",  x"fe",  x"42",  x"c2",  x"04", -- 1EE8
         x"3f",  x"3a",  x"fa",  x"f0",  x"fe",  x"46",  x"c2",  x"4c", -- 1EF0
         x"39",  x"3a",  x"6b",  x"f1",  x"fe",  x"04",  x"da",  x"4c", -- 1EF8
         x"39",  x"c3",  x"0a",  x"3f",  x"79",  x"fe",  x"4a",  x"c2", -- 1F00
         x"4c",  x"39",  x"cd",  x"10",  x"3f",  x"c3",  x"41",  x"3d", -- 1F08
         x"79",  x"32",  x"a6",  x"f1",  x"af",  x"32",  x"13",  x"f1", -- 1F10
         x"c9",  x"3a",  x"0b",  x"f1",  x"d6",  x"31",  x"87",  x"5f", -- 1F18
         x"16",  x"00",  x"21",  x"22",  x"1a",  x"19",  x"5e",  x"23", -- 1F20
         x"56",  x"eb",  x"22",  x"05",  x"f0",  x"cd",  x"03",  x"f0", -- 1F28
         x"c9",  x"cd",  x"36",  x"21",  x"af",  x"32",  x"13",  x"f1", -- 1F30
         x"3e",  x"38",  x"32",  x"0b",  x"f1",  x"32",  x"ec",  x"f0", -- 1F38
         x"21",  x"68",  x"78",  x"22",  x"6b",  x"f1",  x"22",  x"6d", -- 1F40
         x"f1",  x"21",  x"98",  x"98",  x"22",  x"5b",  x"f1",  x"21", -- 1F48
         x"a8",  x"a8",  x"22",  x"5d",  x"f1",  x"21",  x"8e",  x"17", -- 1F50
         x"11",  x"7b",  x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"15", -- 1F58
         x"f1",  x"c3",  x"4c",  x"39",  x"3a",  x"13",  x"f1",  x"b7", -- 1F60
         x"ca",  x"4c",  x"39",  x"c9",  x"3e",  x"3b",  x"32",  x"0b", -- 1F68
         x"f1",  x"32",  x"ec",  x"f0",  x"cd",  x"36",  x"21",  x"cd", -- 1F70
         x"85",  x"21",  x"21",  x"27",  x"37",  x"22",  x"6f",  x"f1", -- 1F78
         x"21",  x"0b",  x"88",  x"22",  x"71",  x"f1",  x"21",  x"d7", -- 1F80
         x"e7",  x"22",  x"74",  x"f1",  x"22",  x"76",  x"f1",  x"22", -- 1F88
         x"78",  x"f1",  x"21",  x"a7",  x"a7",  x"22",  x"5b",  x"f1", -- 1F90
         x"21",  x"b7",  x"b7",  x"22",  x"5d",  x"f1",  x"21",  x"4f", -- 1F98
         x"4f",  x"22",  x"5f",  x"f1",  x"22",  x"68",  x"f1",  x"21", -- 1FA0
         x"4a",  x"80",  x"22",  x"61",  x"f1",  x"21",  x"37",  x"37", -- 1FA8
         x"22",  x"64",  x"f1",  x"21",  x"47",  x"47",  x"22",  x"66", -- 1FB0
         x"f1",  x"cd",  x"a5",  x"21",  x"21",  x"43",  x"63",  x"22", -- 1FB8
         x"7f",  x"f1",  x"22",  x"88",  x"f1",  x"21",  x"74",  x"16", -- 1FC0
         x"11",  x"84",  x"f1",  x"cd",  x"4d",  x"1b",  x"3e",  x"1f", -- 1FC8
         x"32",  x"81",  x"f1",  x"21",  x"09",  x"09",  x"22",  x"92", -- 1FD0
         x"f1",  x"22",  x"94",  x"f1",  x"22",  x"96",  x"f1",  x"21", -- 1FD8
         x"ca",  x"44",  x"22",  x"17",  x"f1",  x"3e",  x"01",  x"32", -- 1FE0
         x"1a",  x"f1",  x"01",  x"9c",  x"f1",  x"21",  x"a2",  x"f1", -- 1FE8
         x"cd",  x"6d",  x"12",  x"af",  x"32",  x"e8",  x"f0",  x"cd", -- 1FF0
         x"42",  x"44",  x"cd",  x"9f",  x"1a",  x"c3",  x"4c",  x"39"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
