library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_a5 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_a5;

architecture rtl of rom_a5 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0000
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0010
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0028
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0038
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0048
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0050
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0068
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0078
         x"ff",  x"fe",  x"fe",  x"ff",  x"ff",  x"ff",  x"fe",  x"fe", -- 0080
         x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"ff",  x"ff",  x"fe", -- 0088
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0090
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0098
         x"ff",  x"ff",  x"ef",  x"f7",  x"fb",  x"fd",  x"fe",  x"fe", -- 00A0
         x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00A8
         x"ff",  x"ff",  x"ef",  x"f7",  x"fb",  x"fd",  x"fc",  x"fc", -- 00B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fc",  x"ff", -- 00C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"e4",  x"e4",  x"e4",  x"ff", -- 00E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00E8
         x"ff",  x"ff",  x"ff",  x"eb",  x"c3",  x"f3",  x"ff",  x"ff", -- 00F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 00F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0100
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0108
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0110
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0130
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0140
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0148
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0150
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0160
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0170
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0178
         x"c0",  x"c0",  x"ff",  x"fe",  x"fe",  x"fe",  x"fd",  x"fc", -- 0180
         x"fe",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"fd",  x"fd", -- 0188
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f7",  x"f7",  x"e1", -- 0190
         x"07",  x"17",  x"1f",  x"3c",  x"00",  x"80",  x"fc",  x"ff", -- 0198
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f8",  x"f8", -- 01A0
         x"f0",  x"f9",  x"c1",  x"f0",  x"ff",  x"f8",  x"ff",  x"ff", -- 01A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"f8", -- 01B0
         x"ff",  x"c0",  x"e7",  x"ff",  x"ff",  x"f0",  x"ff",  x"ff", -- 01B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01C8
         x"ff",  x"ff",  x"ff",  x"f5",  x"e1",  x"f9",  x"ff",  x"ff", -- 01D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01D8
         x"ff",  x"f3",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 01E0
         x"00",  x"00",  x"00",  x"00",  x"80",  x"80",  x"c0",  x"c1", -- 01E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0200
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0210
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0220
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0230
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0238
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0240
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0268
         x"e4",  x"e5",  x"e7",  x"e7",  x"ff",  x"ff",  x"ff",  x"ff", -- 0270
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0278
         x"00",  x"00",  x"fd",  x"f0",  x"ca",  x"81",  x"44",  x"be", -- 0280
         x"be",  x"35",  x"7f",  x"ff",  x"ff",  x"ef",  x"ff",  x"ff", -- 0288
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0290
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0298
         x"ff",  x"ff",  x"ff",  x"ff",  x"df",  x"ec",  x"e4",  x"f0", -- 02A0
         x"f0",  x"f9",  x"ff",  x"ff",  x"fe",  x"fd",  x"ff",  x"ff", -- 02A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"f1",  x"f1",  x"21",  x"31", -- 02B0
         x"c1",  x"fd",  x"c1",  x"e7",  x"fe",  x"fd",  x"ff",  x"ff", -- 02B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"fa",  x"f0",  x"fc",  x"ff", -- 02C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02C8
         x"ff",  x"f3",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 02D0
         x"92",  x"92",  x"fe",  x"7c",  x"fc",  x"b8",  x"c0",  x"c1", -- 02D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0300
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0308
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0310
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0318
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0320
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0328
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0330
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0338
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0340
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0348
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0350
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0358
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0360
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0368
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0370
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0378
         x"c0",  x"c0",  x"ff",  x"ff",  x"ff",  x"fc",  x"fd",  x"fe", -- 0380
         x"fe",  x"fe",  x"fc",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0388
         x"7e",  x"1e",  x"0c",  x"c0",  x"c0",  x"00",  x"03",  x"3f", -- 0390
         x"1f",  x"3f",  x"3f",  x"7f",  x"7f",  x"ff",  x"ff",  x"7f", -- 0398
         x"ff",  x"ff",  x"ef",  x"f7",  x"fb",  x"fd",  x"fc",  x"fc", -- 03A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"fe", -- 03B0
         x"fe",  x"fe",  x"fd",  x"e3",  x"f3",  x"ff",  x"ff",  x"ff", -- 03B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"3f",  x"0f",  x"07", -- 03C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fd",  x"f8",  x"fe", -- 03E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0400
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0408
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0410
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0418
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0420
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0428
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0430
         x"ff",  x"f8",  x"f8",  x"f8",  x"f8",  x"f8",  x"f8",  x"ff", -- 0438
         x"ff",  x"ff",  x"ff",  x"ff",  x"e0",  x"ff",  x"ff",  x"ff", -- 0440
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0448
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0450
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0458
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"f0",  x"e4", -- 0460
         x"ee",  x"e7",  x"e7",  x"e6",  x"f0",  x"f9",  x"ff",  x"ff", -- 0468
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0470
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f7", -- 0478
         x"00",  x"00",  x"f1",  x"ca",  x"e1",  x"f1",  x"b5",  x"77", -- 0480
         x"1f",  x"df",  x"ff",  x"7f",  x"df",  x"fd",  x"f7",  x"ff", -- 0488
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0490
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f0",  x"e9",  x"c4", -- 0498
         x"ff",  x"1f",  x"ff",  x"ff",  x"fc",  x"ff",  x"ff",  x"ff", -- 04A0
         x"fe",  x"fd",  x"f3",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 04A8
         x"f8",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fb",  x"fb", -- 04B0
         x"ff",  x"fd",  x"f3",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 04B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"df",  x"cf",  x"c3",  x"81", -- 04C0
         x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"01", -- 04C8
         x"03",  x"01",  x"00",  x"00",  x"00",  x"80",  x"c0",  x"e0", -- 04D0
         x"e0",  x"f0",  x"f8",  x"fc",  x"fe",  x"ff",  x"ff",  x"ff", -- 04D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"01",  x"c0",  x"81",  x"c0", -- 04E0
         x"62",  x"00",  x"87",  x"bf",  x"ff",  x"ff",  x"ff",  x"ff", -- 04E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"c0", -- 04F0
         x"62",  x"00",  x"87",  x"bf",  x"ff",  x"ff",  x"ff",  x"ff", -- 04F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0500
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0508
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0510
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0518
         x"ff",  x"fe",  x"fc",  x"fc",  x"fc",  x"fc",  x"ff",  x"ff", -- 0520
         x"f3",  x"f7",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0528
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0530
         x"ff",  x"ff",  x"7f",  x"1f",  x"97",  x"01",  x"47",  x"8c", -- 0538
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0540
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0548
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0550
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0558
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0560
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0568
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0570
         x"ff",  x"ff",  x"ff",  x"f7",  x"f3",  x"f9",  x"fc",  x"e0", -- 0578
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0580
         x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"ff",  x"ff",  x"fe", -- 0588
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc", -- 0590
         x"f8",  x"f8",  x"f8",  x"fc",  x"f0",  x"f1",  x"cb",  x"e7", -- 0598
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7c", -- 05A0
         x"06",  x"80",  x"a1",  x"c0",  x"00",  x"ff",  x"ff",  x"ff", -- 05A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7c", -- 05B0
         x"06",  x"80",  x"a3",  x"c3",  x"81",  x"c0",  x"01",  x"ff", -- 05B8
         x"ff",  x"f3",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 05C0
         x"00",  x"4e",  x"ff",  x"ff",  x"ff",  x"f8",  x"f8",  x"c1", -- 05C8
         x"ff",  x"f0",  x"e0",  x"f0",  x"c0",  x"e0",  x"e0",  x"e0", -- 05D0
         x"c0",  x"e0",  x"f0",  x"fc",  x"f8",  x"fd",  x"fb",  x"ff", -- 05D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc",  x"fe",  x"fe", -- 05E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 05E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 05F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 05F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0600
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0608
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0610
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0618
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0620
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0628
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0630
         x"ff",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88",  x"ff", -- 0638
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0640
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0648
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0650
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"80",  x"00",  x"ff", -- 0658
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0660
         x"ff",  x"ff",  x"3f",  x"5f",  x"1f",  x"47",  x"1f",  x"23", -- 0668
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0670
         x"fe",  x"ff",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0678
         x"ff",  x"d7",  x"c7",  x"d1",  x"80",  x"c1",  x"91",  x"b0", -- 0680
         x"a4",  x"6f",  x"63",  x"c7",  x"c3",  x"48",  x"54",  x"83", -- 0688
         x"cf",  x"8f",  x"c4",  x"e0",  x"f8",  x"7c",  x"3c",  x"10", -- 0690
         x"06",  x"0f",  x"00",  x"f0",  x"f9",  x"fc",  x"ff",  x"ff", -- 0698
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc",  x"f8", -- 06A0
         x"f8",  x"f8",  x"fc",  x"fc",  x"f8",  x"fa",  x"fc",  x"fe", -- 06A8
         x"7f",  x"bf",  x"8f",  x"07",  x"03",  x"81",  x"f1",  x"fb", -- 06B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 06B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc",  x"f8", -- 06C0
         x"f8",  x"f8",  x"fc",  x"fc",  x"f8",  x"fa",  x"fc",  x"fe", -- 06C8
         x"bf",  x"bf",  x"8f",  x"0f",  x"07",  x"07",  x"83",  x"e3", -- 06D0
         x"eb",  x"ff",  x"ff",  x"3f",  x"bf",  x"7f",  x"ff",  x"ff", -- 06D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 06E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 06E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 06F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 06F8
         x"ff",  x"fe",  x"fc",  x"fc",  x"fc",  x"fc",  x"ff",  x"df", -- 0700
         x"ef",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0708
         x"ff",  x"ff",  x"7e",  x"7e",  x"7e",  x"fe",  x"fc",  x"fd", -- 0710
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0718
         x"ff",  x"ff",  x"f9",  x"f7",  x"fe",  x"fc",  x"f1",  x"fb", -- 0720
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0728
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0730
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0738
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0740
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0748
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0750
         x"ff",  x"ff",  x"ff",  x"ff",  x"fd",  x"00",  x"00",  x"ff", -- 0758
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0760
         x"ff",  x"ff",  x"c7",  x"c7",  x"c3",  x"e3",  x"f3",  x"ff", -- 0768
         x"23",  x"01",  x"01",  x"00",  x"00",  x"00",  x"00",  x"06", -- 0770
         x"0f",  x"0f",  x"0f",  x"0f",  x"07",  x"03",  x"03",  x"0f", -- 0778
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fc", -- 0780
         x"e4",  x"f0",  x"f9",  x"f3",  x"ff",  x"ff",  x"ff",  x"ff", -- 0788
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0790
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0798
         x"4f",  x"06",  x"00",  x"87",  x"cf",  x"ff",  x"ff",  x"ff", -- 07A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"f7",  x"f3",  x"f8",  x"fc", -- 07B8
         x"ff",  x"ff",  x"ff",  x"fa",  x"f0",  x"fc",  x"ff",  x"ff", -- 07C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 07E8
         x"04",  x"00",  x"00",  x"00",  x"01",  x"01",  x"04",  x"06", -- 07F0
         x"0f",  x"0b",  x"03",  x"07",  x"07",  x"03",  x"03",  x"0f", -- 07F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f", -- 0800
         x"1f",  x"1f",  x"7f",  x"7f",  x"ff",  x"7f",  x"3f",  x"3f", -- 0808
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0810
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0818
         x"1f",  x"3f",  x"1f",  x"3f",  x"1f",  x"1f",  x"3f",  x"1f", -- 0820
         x"3f",  x"3f",  x"1f",  x"3f",  x"3f",  x"3f",  x"ff",  x"ff", -- 0828
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0830
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0838
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0840
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0848
         x"83",  x"c7",  x"ef",  x"cf",  x"ef",  x"ff",  x"ff",  x"bf", -- 0850
         x"bf",  x"ff",  x"ff",  x"ff",  x"ef",  x"cf",  x"ff",  x"ff", -- 0858
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0860
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0868
         x"00",  x"f8",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"3f", -- 0870
         x"1f",  x"1f",  x"bf",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0878
         x"ff",  x"ff",  x"ff",  x"ff",  x"f7",  x"f7",  x"e1",  x"03", -- 0880
         x"10",  x"78",  x"0c",  x"1f",  x"9f",  x"9f",  x"ff",  x"ff", -- 0888
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe", -- 0890
         x"fe",  x"fc",  x"e0",  x"e2",  x"f1",  x"f3",  x"f3",  x"f1", -- 0898
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f", -- 0900
         x"1f",  x"1f",  x"7f",  x"7f",  x"ff",  x"7f",  x"3f",  x"00", -- 0908
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0910
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0918
         x"00",  x"01",  x"01",  x"3f",  x"1f",  x"1f",  x"3f",  x"1f", -- 0920
         x"3f",  x"3f",  x"1f",  x"3f",  x"3f",  x"3f",  x"ff",  x"ff", -- 0928
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc",  x"f8", -- 0930
         x"f8",  x"f0",  x"f0",  x"f0",  x"f0",  x"f8",  x"f8",  x"ff", -- 0938
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0940
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fc", -- 0948
         x"f9",  x"f3",  x"f2",  x"f8",  x"fc",  x"ff",  x"fc",  x"f8", -- 0950
         x"f8",  x"f8",  x"f4",  x"f0",  x"d0",  x"cb",  x"fd",  x"fe", -- 0958
         x"f9",  x"7c",  x"38",  x"20",  x"04",  x"0f",  x"0f",  x"0f", -- 0960
         x"0f",  x"1d",  x"dd",  x"b1",  x"bf",  x"7f",  x"ff",  x"7f", -- 0968
         x"c0",  x"c0",  x"ff",  x"fe",  x"fd",  x"fe",  x"ff",  x"fe", -- 0970
         x"fe",  x"fd",  x"fd",  x"fd",  x"fd",  x"fd",  x"fd",  x"ff", -- 0978
         x"ff",  x"ff",  x"dd",  x"c4",  x"f4",  x"f0",  x"f9",  x"ff", -- 0980
         x"fe",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0988
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0990
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0998
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 09F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A00
         x"f7",  x"f7",  x"eb",  x"ff",  x"eb",  x"c1",  x"80",  x"80", -- 0A08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0A20
         x"00",  x"00",  x"41",  x"c1",  x"c1",  x"c1",  x"80",  x"00", -- 0A28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A38
         x"f9",  x"f3",  x"f2",  x"f8",  x"fc",  x"ff",  x"fc",  x"f8", -- 0A40
         x"f8",  x"f8",  x"f4",  x"f0",  x"d0",  x"cb",  x"fd",  x"fe", -- 0A48
         x"ff",  x"1f",  x"3f",  x"3f",  x"8f",  x"07",  x"03",  x"91", -- 0A50
         x"f1",  x"7b",  x"7f",  x"ff",  x"7f",  x"ff",  x"ff",  x"ff", -- 0A58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A60
         x"ff",  x"ff",  x"ff",  x"fa",  x"f0",  x"e0",  x"e0",  x"f0", -- 0A68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A70
         x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"e0",  x"e0", -- 0A78
         x"ff",  x"ff",  x"ff",  x"ff",  x"f7",  x"f7",  x"e1",  x"07", -- 0A80
         x"1f",  x"7f",  x"3f",  x"bf",  x"7f",  x"ff",  x"ff",  x"ff", -- 0A88
         x"f8",  x"1c",  x"0f",  x"0f",  x"00",  x"00",  x"00",  x"c0", -- 0A90
         x"e0",  x"e0",  x"f8",  x"fc",  x"ff",  x"ff",  x"ff",  x"ff", -- 0A98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0AF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B38
         x"ff",  x"1f",  x"3f",  x"3f",  x"8f",  x"07",  x"03",  x"91", -- 0B40
         x"f1",  x"7b",  x"7f",  x"ff",  x"7f",  x"ff",  x"ff",  x"ff", -- 0B48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B60
         x"ff",  x"ef",  x"ef",  x"c3",  x"0f",  x"0f",  x"07",  x"d7", -- 0B68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B70
         x"ff",  x"ff",  x"7f",  x"1f",  x"97",  x"01",  x"47",  x"84", -- 0B78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B80
         x"ff",  x"ff",  x"ff",  x"ff",  x"fb",  x"fd",  x"f0",  x"fc", -- 0B88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C30
         x"ff",  x"f7",  x"e3",  x"e7",  x"c1",  x"c1",  x"9c",  x"a2", -- 0C38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C50
         x"bf",  x"8f",  x"3f",  x"3f",  x"ff",  x"7f",  x"ff",  x"6f", -- 0C58
         x"fd",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C68
         x"04",  x"04",  x"09",  x"00",  x"00",  x"00",  x"03",  x"0e", -- 0C70
         x"0f",  x"0f",  x"0f",  x"0f",  x"07",  x"03",  x"03",  x"0f", -- 0C78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C80
         x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"fc",  x"e0",  x"e0", -- 0C88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fd", -- 0C98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"df",  x"c7",  x"9f", -- 0D40
         x"1f",  x"7f",  x"3f",  x"3f",  x"bf",  x"b7",  x"80",  x"81", -- 0D48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe", -- 0D50
         x"fc",  x"f8",  x"f0",  x"f1",  x"f3",  x"ff",  x"ff",  x"ff", -- 0D58
         x"6f",  x"7f",  x"7f",  x"fb",  x"e3",  x"e1",  x"c0",  x"80", -- 0D60
         x"80",  x"80",  x"c1",  x"e1",  x"f1",  x"c7",  x"e3",  x"f8", -- 0D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D80
         x"ff",  x"ff",  x"ff",  x"f8",  x"f8",  x"fc",  x"fc",  x"fc", -- 0D88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"e3",  x"c1",  x"c0", -- 0D90
         x"c4",  x"e4",  x"ec",  x"fb",  x"f3",  x"f3",  x"f9",  x"fc", -- 0D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E28
         x"22",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E30
         x"00",  x"41",  x"00",  x"41",  x"c1",  x"d5",  x"94",  x"36", -- 0E38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E48
         x"77",  x"71",  x"70",  x"f0",  x"60",  x"27",  x"03",  x"01", -- 0E50
         x"00",  x"00",  x"31",  x"38",  x"3e",  x"fe",  x"7d",  x"1c", -- 0E58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E60
         x"ff",  x"ff",  x"df",  x"c7",  x"9f",  x"9f",  x"7c",  x"00", -- 0E68
         x"10",  x"21",  x"01",  x"01",  x"07",  x"09",  x"04",  x"0e", -- 0E70
         x"0f",  x"0f",  x"0f",  x"0f",  x"07",  x"03",  x"03",  x"0f", -- 0E78
         x"fc",  x"fe",  x"fe",  x"ff",  x"ff",  x"fe",  x"fc",  x"f8", -- 0E80
         x"f8",  x"f8",  x"f8",  x"fc",  x"fe",  x"f8",  x"fc",  x"fe", -- 0E88
         x"7d",  x"78",  x"01",  x"89",  x"ef",  x"1f",  x"3f",  x"1f", -- 0E90
         x"0f",  x"07",  x"c7",  x"ef",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0EF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F08
         x"ff",  x"ff",  x"ff",  x"f5",  x"e1",  x"f9",  x"ff",  x"ff", -- 0F10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F38
         x"f9",  x"7c",  x"38",  x"20",  x"04",  x"0f",  x"0f",  x"0f", -- 0F40
         x"0f",  x"1d",  x"dd",  x"b1",  x"bf",  x"7f",  x"ff",  x"7f", -- 0F48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F58
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"c6",  x"82",  x"82", -- 0F60
         x"86",  x"cc",  x"cc",  x"ee",  x"e7",  x"e7",  x"f3",  x"f8", -- 0F68
         x"00",  x"00",  x"fd",  x"f0",  x"88",  x"a5",  x"54",  x"b7", -- 0F70
         x"3f",  x"ff",  x"df",  x"ff",  x"f7",  x"ff",  x"fb",  x"ff", -- 0F78
         x"ff",  x"ff",  x"3f",  x"1f",  x"bf",  x"ff",  x"ff",  x"ff", -- 0F80
         x"7f",  x"7f",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f",  x"9f", -- 0F88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc", -- 0F90
         x"fc",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1000
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1010
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1028
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1038
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1048
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1050
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1068
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1078
         x"7f",  x"7f",  x"ff",  x"7f",  x"ff",  x"ff",  x"ff",  x"7f", -- 1080
         x"7f",  x"7f",  x"ff",  x"7f",  x"ff",  x"7f",  x"7f",  x"ff", -- 1088
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1090
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1098
         x"ff",  x"ff",  x"ff",  x"ff",  x"c7",  x"c7",  x"87",  x"47", -- 10A0
         x"0f",  x"9d",  x"ff",  x"83",  x"fb",  x"fb",  x"ff",  x"ff", -- 10A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"8f",  x"8f",  x"0f",  x"1f", -- 10B0
         x"3b",  x"fb",  x"bf",  x"ff",  x"c3",  x"bf",  x"ff",  x"ff", -- 10B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"bf",  x"3f",  x"3f", -- 10C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 10D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"27",  x"27", -- 10D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ea", -- 10E0
         x"c2",  x"f2",  x"ff",  x"fe",  x"fe",  x"fe",  x"ff",  x"fa", -- 10E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ae", -- 10F0
         x"0f",  x"cf",  x"ff",  x"ff",  x"fe",  x"fe",  x"ff",  x"fa", -- 10F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1100
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1108
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1110
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1128
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1130
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1138
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1140
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1148
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1150
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1160
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1170
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1178
         x"00",  x"00",  x"cf",  x"0f",  x"e3",  x"8b",  x"15",  x"f8", -- 1180
         x"7c",  x"fe",  x"df",  x"ff",  x"ff",  x"fe",  x"fa",  x"ff", -- 1188
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1190
         x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"0f",  x"01", -- 1198
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 11A0
         x"ff",  x"ff",  x"43",  x"7f",  x"ff",  x"03",  x"ff",  x"ff", -- 11A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"1f",  x"1f",  x"19",  x"00", -- 11B0
         x"63",  x"7f",  x"ff",  x"ff",  x"ff",  x"1f",  x"ff",  x"ff", -- 11B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 11C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 11C8
         x"27",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe", -- 11D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"ff",  x"fa", -- 11D8
         x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f",  x"3f",  x"1f", -- 11E0
         x"0f",  x"0f",  x"0f",  x"0f",  x"27",  x"27",  x"37",  x"57", -- 11E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 11F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 11F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1200
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1210
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1220
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1230
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1238
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1240
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1268
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1270
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1278
         x"03",  x"03",  x"ff",  x"7f",  x"7f",  x"3f",  x"7f",  x"7f", -- 1280
         x"3f",  x"bf",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1288
         x"fc",  x"fc",  x"fe",  x"ff",  x"ff",  x"ff",  x"fe",  x"fc", -- 1290
         x"fc",  x"fc",  x"fe",  x"fe",  x"fe",  x"fc",  x"fc",  x"fc", -- 1298
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f", -- 12A0
         x"df",  x"df",  x"f7",  x"ef",  x"1f",  x"ff",  x"ff",  x"ff", -- 12A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 12B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"1f",  x"e7",  x"ff",  x"ff", -- 12B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe", -- 12C0
         x"fe",  x"fc",  x"7f",  x"ff",  x"fe",  x"fe",  x"ff",  x"fa", -- 12C8
         x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f",  x"3f",  x"1f", -- 12D0
         x"0f",  x"0f",  x"0f",  x"0f",  x"27",  x"27",  x"37",  x"57", -- 12D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 12E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 12E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 12F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 12F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1300
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1308
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1310
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1318
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1320
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1328
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1330
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1338
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1340
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1348
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1350
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1358
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1360
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1368
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1370
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1378
         x"00",  x"00",  x"9f",  x"cb",  x"3f",  x"47",  x"0d",  x"3b", -- 1380
         x"bb",  x"ff",  x"fe",  x"be",  x"be",  x"ee",  x"ff",  x"7e", -- 1388
         x"00",  x"80",  x"fd",  x"bf",  x"5f",  x"1f",  x"df",  x"9f", -- 1390
         x"1f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1398
         x"ff",  x"ff",  x"ff",  x"ff",  x"8f",  x"8f",  x"0f",  x"1f", -- 13A0
         x"3f",  x"ff",  x"9f",  x"ef",  x"c3",  x"bf",  x"ff",  x"ff", -- 13A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"3f",  x"3f",  x"3f",  x"3f", -- 13B0
         x"bf",  x"df",  x"ef",  x"27",  x"27",  x"2f",  x"ff",  x"ff", -- 13B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 13C0
         x"ff",  x"ff",  x"fe",  x"e0",  x"f0",  x"f8",  x"fe",  x"ff", -- 13C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 13D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"af",  x"0f",  x"cf", -- 13D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 13E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f", -- 13E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 13F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 13F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1400
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1408
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1410
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1418
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 1420
         x"bf",  x"ff",  x"fb",  x"fb",  x"ff",  x"ff",  x"ff",  x"ff", -- 1428
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1430
         x"ff",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88",  x"ff", -- 1438
         x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"ff",  x"ff",  x"ff", -- 1440
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1448
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1450
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1458
         x"ff",  x"ff",  x"bf",  x"7f",  x"ff",  x"ff",  x"ff",  x"7f", -- 1460
         x"7f",  x"7f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1468
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1470
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1478
         x"03",  x"03",  x"ff",  x"7f",  x"3f",  x"bf",  x"3f",  x"ff", -- 1480
         x"ff",  x"bf",  x"ff",  x"bf",  x"3f",  x"ff",  x"ff",  x"ff", -- 1488
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1490
         x"ff",  x"ff",  x"bf",  x"bf",  x"0f",  x"3f",  x"ff",  x"ff", -- 1498
         x"ff",  x"ff",  x"ff",  x"df",  x"3f",  x"7f",  x"ff",  x"ff", -- 14A0
         x"3f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 14A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"bf", -- 14B0
         x"bf",  x"df",  x"df",  x"df",  x"ff",  x"ff",  x"ff",  x"ff", -- 14B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 14C0
         x"7f",  x"1f",  x"1f",  x"1f",  x"3f",  x"7f",  x"ff",  x"ff", -- 14C8
         x"ff",  x"ff",  x"ff",  x"3f",  x"79",  x"ff",  x"f9",  x"d0", -- 14D0
         x"d0",  x"f9",  x"ff",  x"f9",  x"7f",  x"3f",  x"ff",  x"ff", -- 14D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f7", -- 14E0
         x"c1",  x"05",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 14E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f7", -- 14F0
         x"c1",  x"05",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 14F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1500
         x"e7",  x"d5",  x"d8",  x"fe",  x"fc",  x"fe",  x"ff",  x"ff", -- 1508
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1510
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1518
         x"ff",  x"ff",  x"9f",  x"bf",  x"ff",  x"fd",  x"ff",  x"ff", -- 1520
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1528
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1530
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 1538
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1540
         x"df",  x"f7",  x"bd",  x"ef",  x"c7",  x"ef",  x"ef",  x"ef", -- 1548
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1550
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1558
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1560
         x"fd",  x"fc",  x"fe",  x"fe",  x"fe",  x"ff",  x"ff",  x"ff", -- 1568
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1570
         x"ff",  x"ff",  x"ff",  x"cf",  x"8f",  x"0f",  x"0f",  x"01", -- 1578
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1580
         x"7f",  x"7f",  x"ff",  x"7f",  x"ff",  x"7f",  x"7f",  x"ff", -- 1588
         x"ff",  x"ff",  x"ff",  x"fd",  x"fc",  x"f8",  x"f8",  x"60", -- 1590
         x"00",  x"00",  x"00",  x"3d",  x"7f",  x"ff",  x"ff",  x"ff", -- 1598
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f7", -- 15A0
         x"c1",  x"05",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f7", -- 15B0
         x"c1",  x"05",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15B8
         x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"7f",  x"3f",  x"1f", -- 15C0
         x"0f",  x"0f",  x"0f",  x"0f",  x"27",  x"27",  x"37",  x"57", -- 15C8
         x"ff",  x"5f",  x"37",  x"0f",  x"0f",  x"0f",  x"07",  x"0f", -- 15D0
         x"07",  x"07",  x"0f",  x"0f",  x"8f",  x"0f",  x"1f",  x"3f", -- 15D8
         x"3f",  x"3f",  x"7f",  x"7f",  x"7f",  x"7f",  x"7f",  x"3f", -- 15E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ef",  x"ef", -- 1600
         x"df",  x"ff",  x"fb",  x"fb",  x"ff",  x"ff",  x"ff",  x"ff", -- 1608
         x"ff",  x"fc",  x"f3",  x"ff",  x"ff",  x"ff",  x"3f",  x"df", -- 1610
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1618
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc",  x"ff",  x"ff", -- 1620
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1628
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1630
         x"ff",  x"8f",  x"8f",  x"8f",  x"8f",  x"8f",  x"8f",  x"ff", -- 1638
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1640
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1648
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1650
         x"ff",  x"ff",  x"ff",  x"ff",  x"fd",  x"00",  x"00",  x"ff", -- 1658
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1660
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1668
         x"fe",  x"fe",  x"fc",  x"f8",  x"d0",  x"c0",  x"80",  x"00", -- 1670
         x"82",  x"4e",  x"ae",  x"6e",  x"fe",  x"fc",  x"f8",  x"e0", -- 1678
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1680
         x"ff",  x"ff",  x"ff",  x"bf",  x"7f",  x"1d",  x"01",  x"00", -- 1688
         x"ff",  x"ff",  x"ff",  x"7f",  x"ff",  x"3f",  x"1f",  x"0f", -- 1690
         x"07",  x"c7",  x"6f",  x"7f",  x"7f",  x"ff",  x"ff",  x"ff", -- 1698
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fc",  x"40",  x"00", -- 16A0
         x"00",  x"00",  x"38",  x"3c",  x"7c",  x"fc",  x"fc",  x"3c", -- 16A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fc",  x"40",  x"00", -- 16C0
         x"00",  x"00",  x"38",  x"3d",  x"7d",  x"fd",  x"fd",  x"3c", -- 16C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fb",  x"fb",  x"f0", -- 16E0
         x"83",  x"cf",  x"c7",  x"ff",  x"e7",  x"e3",  x"e1",  x"f0", -- 16E8
         x"f8",  x"fc",  x"fe",  x"fc",  x"f9",  x"c1",  x"c3",  x"e3", -- 16F0
         x"e3",  x"e3",  x"e7",  x"e7",  x"e7",  x"ef",  x"ff",  x"ff", -- 16F8
         x"ff",  x"ff",  x"9f",  x"bf",  x"ff",  x"fd",  x"ff",  x"ff", -- 1700
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1708
         x"ff",  x"7f",  x"4f",  x"5f",  x"7f",  x"7e",  x"ff",  x"7f", -- 1710
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1718
         x"ff",  x"7f",  x"8f",  x"df",  x"df",  x"be",  x"bf",  x"bf", -- 1720
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1728
         x"fe",  x"fe",  x"fc",  x"fc",  x"fc",  x"fc",  x"fc",  x"fe", -- 1730
         x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fc",  x"f8",  x"e0", -- 1738
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1740
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1748
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1750
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"07",  x"03",  x"ff", -- 1758
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1760
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1768
         x"ff",  x"ff",  x"ff",  x"df",  x"1f",  x"0f",  x"07",  x"0b", -- 1770
         x"97",  x"ab",  x"b7",  x"ff",  x"ff",  x"ff",  x"bf",  x"7f", -- 1778
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"79",  x"79",  x"78", -- 1780
         x"79",  x"f8",  x"fc",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1788
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1790
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1798
         x"3f",  x"7f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"cf",  x"0f",  x"0f", -- 17B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ea", -- 17C0
         x"c2",  x"f2",  x"ff",  x"fe",  x"fe",  x"fe",  x"ff",  x"fa", -- 17C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17D8
         x"fe",  x"fe",  x"fc",  x"fc",  x"fc",  x"fc",  x"fc",  x"fc", -- 17E0
         x"fe",  x"fe",  x"fe",  x"fe",  x"fe",  x"fc",  x"f8",  x"e0", -- 17E8
         x"3f",  x"3f",  x"3f",  x"7f",  x"ff",  x"7f",  x"7f",  x"7f", -- 17F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"bf",  x"7f", -- 17F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1800
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1808
         x"e0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"c0", -- 1810
         x"c0",  x"c0",  x"80",  x"c4",  x"ec",  x"fc",  x"ff",  x"fe", -- 1818
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1820
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1828
         x"ff",  x"ff",  x"ff",  x"ff",  x"e0",  x"c0",  x"c0",  x"c0", -- 1830
         x"e0",  x"f0",  x"fc",  x"f9",  x"f9",  x"f8",  x"e0",  x"e0", -- 1838
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1840
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1848
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1850
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1858
         x"80",  x"c0",  x"f8",  x"fc",  x"ff",  x"f0",  x"c0",  x"80", -- 1860
         x"80",  x"82",  x"c7",  x"8f",  x"c3",  x"b9",  x"7e",  x"3e", -- 1868
         x"7f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1870
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1878
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1880
         x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1888
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1890
         x"ff",  x"3f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1898
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1900
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"bf",  x"01", -- 1908
         x"e0",  x"f0",  x"f0",  x"f0",  x"f8",  x"f8",  x"f8",  x"f8", -- 1910
         x"f8",  x"f8",  x"fc",  x"fc",  x"fc",  x"f8",  x"fb",  x"f6", -- 1918
         x"07",  x"af",  x"df",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1920
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1928
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"1f",  x"07", -- 1930
         x"01",  x"00",  x"00",  x"00",  x"00",  x"01",  x"01",  x"03", -- 1938
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1940
         x"fb",  x"f8",  x"f3",  x"83",  x"8f",  x"87",  x"c7",  x"d7", -- 1948
         x"d6",  x"f0",  x"f0",  x"1f",  x"0f",  x"07",  x"02",  x"00", -- 1950
         x"00",  x"00",  x"79",  x"7c",  x"f9",  x"f8",  x"fd",  x"7c", -- 1958
         x"ff",  x"7f",  x"3f",  x"1f",  x"0f",  x"8f",  x"df",  x"ff", -- 1960
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1968
         x"00",  x"00",  x"bf",  x"07",  x"29",  x"55",  x"62",  x"ba", -- 1970
         x"bd",  x"be",  x"fe",  x"fb",  x"ff",  x"ef",  x"ff",  x"ff", -- 1978
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f9",  x"f9",  x"32", -- 1980
         x"66",  x"0e",  x"7f",  x"fd",  x"f8",  x"fc",  x"ff",  x"ff", -- 1988
         x"ff",  x"ff",  x"fe",  x"fe",  x"fa",  x"f8",  x"f8",  x"f9", -- 1990
         x"f9",  x"e3",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1998
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 19F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A08
         x"ff",  x"fe",  x"fe",  x"fc",  x"fc",  x"fc",  x"fc",  x"fc", -- 1A10
         x"fc",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A18
         x"7f",  x"3f",  x"3f",  x"1f",  x"1f",  x"1f",  x"1f",  x"1f", -- 1A20
         x"1f",  x"3f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 1A28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fb",  x"fb",  x"f0", -- 1A30
         x"83",  x"cf",  x"c7",  x"ff",  x"cf",  x"cf",  x"cf",  x"cf", -- 1A38
         x"d6",  x"f0",  x"f0",  x"1f",  x"0f",  x"07",  x"02",  x"00", -- 1A40
         x"00",  x"00",  x"78",  x"7c",  x"f9",  x"f8",  x"fd",  x"7c", -- 1A48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A60
         x"ff",  x"ff",  x"ff",  x"ff",  x"bb",  x"30",  x"20",  x"a0", -- 1A68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A70
         x"ff",  x"ff",  x"ff",  x"bf",  x"8f",  x"01",  x"00",  x"00", -- 1A78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A88
         x"1f",  x"0f",  x"0f",  x"9f",  x"47",  x"03",  x"01",  x"00", -- 1A90
         x"c8",  x"dd",  x"5f",  x"7f",  x"3f",  x"9f",  x"cf",  x"c7", -- 1A98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B28
         x"8f",  x"cf",  x"cf",  x"cf",  x"87",  x"87",  x"87",  x"8f", -- 1B30
         x"8f",  x"8f",  x"9f",  x"9f",  x"9f",  x"df",  x"ff",  x"ff", -- 1B38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B50
         x"ff",  x"ff",  x"ff",  x"f8",  x"f9",  x"f8",  x"f4",  x"c5", -- 1B58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 1B68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 1B78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"cf",  x"0f",  x"0f", -- 1B88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C40
         x"fc",  x"fc",  x"fc",  x"f6",  x"e6",  x"ce",  x"cf",  x"97", -- 1C48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C58
         x"f0",  x"fc",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C68
         x"3f",  x"3f",  x"3f",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f", -- 1C70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"bf",  x"7f", -- 1C78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"3f",  x"87",  x"0f", -- 1C88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D28
         x"ff",  x"fe",  x"fe",  x"fc",  x"fc",  x"fc",  x"fc",  x"fc", -- 1D30
         x"fc",  x"fc",  x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D48
         x"cd",  x"9e",  x"9c",  x"80",  x"80",  x"4c",  x"98",  x"b0", -- 1D50
         x"f0",  x"f0",  x"f8",  x"fc",  x"fe",  x"f8",  x"fc",  x"ff", -- 1D58
         x"bf",  x"8f",  x"81",  x"80",  x"05",  x"3f",  x"1f",  x"0f", -- 1D60
         x"07",  x"07",  x"8f",  x"c7",  x"f3",  x"f3",  x"eb",  x"e4", -- 1D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D80
         x"bf",  x"bf",  x"0f",  x"3f",  x"ff",  x"7f",  x"e7",  x"c3", -- 1D88
         x"fc",  x"f8",  x"f1",  x"f1",  x"18",  x"08",  x"0e",  x"00", -- 1D90
         x"04",  x"06",  x"0f",  x"0f",  x"e7",  x"f7",  x"f3",  x"71", -- 1D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E28
         x"7f",  x"3f",  x"3f",  x"1f",  x"1f",  x"1f",  x"1f",  x"1f", -- 1E30
         x"1f",  x"1f",  x"3f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E38
         x"80",  x"c0",  x"f8",  x"fc",  x"ff",  x"f0",  x"c0",  x"80", -- 1E40
         x"80",  x"82",  x"c7",  x"8f",  x"c3",  x"b9",  x"7e",  x"9e", -- 1E48
         x"ff",  x"ff",  x"3f",  x"1f",  x"bf",  x"ff",  x"ff",  x"ff", -- 1E50
         x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"ff",  x"7f",  x"9f", -- 1E58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"3f", -- 1E68
         x"3f",  x"3f",  x"3f",  x"7f",  x"ff",  x"7f",  x"7f",  x"7f", -- 1E70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"bf",  x"7f", -- 1E78
         x"83",  x"01",  x"70",  x"e0",  x"00",  x"03",  x"01",  x"00", -- 1E80
         x"00",  x"00",  x"01",  x"38",  x"3c",  x"fe",  x"fd",  x"1c", -- 1E88
         x"ff",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"af", -- 1F08
         x"87",  x"9f",  x"ff",  x"fe",  x"fe",  x"7a",  x"bb",  x"ee", -- 1F10
         x"ff",  x"ff",  x"ff",  x"ff",  x"fe",  x"fe",  x"ff",  x"fa", -- 1F18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F28
         x"ff",  x"ff",  x"ff",  x"ff",  x"e0",  x"c0",  x"c0",  x"c0", -- 1F30
         x"e0",  x"f0",  x"fc",  x"f9",  x"f9",  x"f8",  x"f8",  x"e0", -- 1F38
         x"ff",  x"7f",  x"3f",  x"1f",  x"0f",  x"8f",  x"df",  x"ff", -- 1F40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fc",  x"fc",  x"fe", -- 1F58
         x"fe",  x"ff",  x"ff",  x"7d",  x"1b",  x"18",  x"10",  x"00", -- 1F60
         x"08",  x"0f",  x"0f",  x"1f",  x"cf",  x"ef",  x"e7",  x"e3", -- 1F68
         x"03",  x"03",  x"ff",  x"7f",  x"bf",  x"bf",  x"bf",  x"bf", -- 1F70
         x"ff",  x"7f",  x"7f",  x"ff",  x"bf",  x"ff",  x"bf",  x"ff", -- 1F78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"f5",  x"d0",  x"00", -- 1F90
         x"00",  x"d1",  x"fb",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
