library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_g1 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_g1;

architecture rtl of rom_g1 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"f3",  x"c3",  x"0b",  x"00",  x"6d",  x"7a",  x"87",  x"bf", -- 0000
         x"2b",  x"00",  x"5d",  x"31",  x"7e",  x"e0",  x"3e",  x"9a", -- 0008
         x"d3",  x"d3",  x"db",  x"d2",  x"e6",  x"20",  x"c2",  x"38", -- 0010
         x"00",  x"21",  x"00",  x"e0",  x"3e",  x"aa",  x"77",  x"be", -- 0018
         x"c2",  x"1e",  x"00",  x"2f",  x"77",  x"be",  x"c2",  x"24", -- 0020
         x"00",  x"23",  x"7c",  x"fe",  x"00",  x"c2",  x"1c",  x"00", -- 0028
         x"3e",  x"ff",  x"32",  x"cf",  x"e0",  x"cd",  x"08",  x"0e", -- 0030
         x"af",  x"32",  x"cf",  x"e0",  x"cd",  x"53",  x"07",  x"db", -- 0038
         x"d1",  x"e6",  x"80",  x"ca",  x"40",  x"0e",  x"21",  x"2b", -- 0040
         x"0b",  x"cd",  x"1e",  x"04",  x"cd",  x"3b",  x"04",  x"21", -- 0048
         x"8f",  x"e0",  x"01",  x"83",  x"08",  x"1e",  x"40",  x"cd", -- 0050
         x"2f",  x"08",  x"cd",  x"e8",  x"07",  x"1e",  x"01",  x"01", -- 0058
         x"00",  x"c0",  x"cd",  x"65",  x"05",  x"1c",  x"01",  x"00", -- 0060
         x"c8",  x"cd",  x"65",  x"05",  x"1c",  x"01",  x"00",  x"d0", -- 0068
         x"cd",  x"65",  x"05",  x"1c",  x"01",  x"00",  x"d8",  x"cd", -- 0070
         x"65",  x"05",  x"3e",  x"3e",  x"d3",  x"be",  x"cd",  x"3b", -- 0078
         x"04",  x"21",  x"1b",  x"0b",  x"cd",  x"1e",  x"04",  x"01", -- 0080
         x"4b",  x"0b",  x"11",  x"00",  x"05",  x"cd",  x"b2",  x"04", -- 0088
         x"3e",  x"00",  x"d3",  x"bf",  x"01",  x"b0",  x"a0",  x"21", -- 0090
         x"1b",  x"0b",  x"1e",  x"01",  x"cd",  x"10",  x"05",  x"cd", -- 0098
         x"e9",  x"05",  x"01",  x"dc",  x"d0",  x"1e",  x"00",  x"cd", -- 00A0
         x"10",  x"05",  x"cd",  x"3b",  x"04",  x"01",  x"79",  x"0b", -- 00A8
         x"11",  x"01",  x"07",  x"cd",  x"b2",  x"04",  x"cd",  x"e9", -- 00B0
         x"06",  x"cd",  x"3b",  x"04",  x"01",  x"9f",  x"0b",  x"11", -- 00B8
         x"01",  x"02",  x"cd",  x"b2",  x"04",  x"3e",  x"02",  x"d3", -- 00C0
         x"d2",  x"01",  x"b9",  x"0b",  x"11",  x"00",  x"09",  x"cd", -- 00C8
         x"b2",  x"04",  x"cd",  x"51",  x"06",  x"dc",  x"a9",  x"05", -- 00D0
         x"16",  x"09",  x"cd",  x"94",  x"07",  x"cd",  x"e9",  x"05", -- 00D8
         x"cd",  x"e9",  x"05",  x"af",  x"d3",  x"d2",  x"db",  x"d2", -- 00E0
         x"e6",  x"10",  x"c4",  x"a9",  x"05",  x"01",  x"da",  x"0b", -- 00E8
         x"11",  x"02",  x"09",  x"cd",  x"b2",  x"04",  x"cd",  x"12", -- 00F0
         x"06",  x"dc",  x"bc",  x"05",  x"3e",  x"00",  x"d3",  x"d2", -- 00F8
         x"01",  x"ee",  x"0b",  x"11",  x"02",  x"09",  x"cd",  x"b2", -- 0100
         x"04",  x"cd",  x"dc",  x"05",  x"16",  x"09",  x"cd",  x"94", -- 0108
         x"07",  x"01",  x"1a",  x"0c",  x"11",  x"01",  x"09",  x"cd", -- 0110
         x"b2",  x"04",  x"cd",  x"dc",  x"05",  x"11",  x"02",  x"09", -- 0118
         x"cd",  x"96",  x"07",  x"01",  x"3a",  x"0c",  x"11",  x"01", -- 0120
         x"09",  x"cd",  x"b2",  x"04",  x"cd",  x"1e",  x"06",  x"dc", -- 0128
         x"c2",  x"05",  x"3e",  x"04",  x"d3",  x"d2",  x"01",  x"1e", -- 0130
         x"00",  x"cd",  x"df",  x"05",  x"3e",  x"00",  x"d3",  x"d2", -- 0138
         x"01",  x"50",  x"0c",  x"11",  x"01",  x"09",  x"cd",  x"b2", -- 0140
         x"04",  x"cd",  x"dc",  x"05",  x"16",  x"09",  x"cd",  x"94", -- 0148
         x"07",  x"cd",  x"5d",  x"06",  x"dc",  x"c8",  x"05",  x"01", -- 0150
         x"7a",  x"0c",  x"11",  x"02",  x"09",  x"cd",  x"b2",  x"04", -- 0158
         x"21",  x"df",  x"0a",  x"0e",  x"04",  x"e5",  x"c5",  x"5e", -- 0160
         x"23",  x"56",  x"eb",  x"cd",  x"72",  x"06",  x"c1",  x"e1", -- 0168
         x"23",  x"23",  x"0d",  x"c2",  x"65",  x"01",  x"cd",  x"3b", -- 0170
         x"04",  x"01",  x"a2",  x"0c",  x"11",  x"05",  x"10",  x"cd", -- 0178
         x"b2",  x"04",  x"cd",  x"dc",  x"05",  x"cd",  x"3b",  x"04", -- 0180
         x"01",  x"b7",  x"0c",  x"11",  x"01",  x"04",  x"cd",  x"b2", -- 0188
         x"04",  x"cd",  x"9d",  x"07",  x"01",  x"d3",  x"0c",  x"11", -- 0190
         x"01",  x"06",  x"cd",  x"b2",  x"04",  x"21",  x"00",  x"e1", -- 0198
         x"11",  x"ff",  x"ff",  x"cd",  x"65",  x"04",  x"01",  x"ec", -- 01A0
         x"0c",  x"11",  x"01",  x"08",  x"cd",  x"b2",  x"04",  x"cd", -- 01A8
         x"dc",  x"05",  x"cd",  x"3b",  x"04",  x"01",  x"fc",  x"0c", -- 01B0
         x"11",  x"00",  x"07",  x"cd",  x"b2",  x"04",  x"cd",  x"dc", -- 01B8
         x"05",  x"21",  x"2b",  x"0b",  x"cd",  x"1e",  x"04",  x"0e", -- 01C0
         x"ff",  x"21",  x"00",  x"4c",  x"11",  x"00",  x"50",  x"cd", -- 01C8
         x"c8",  x"06",  x"cd",  x"8f",  x"05",  x"cd",  x"de",  x"06", -- 01D0
         x"0e",  x"10",  x"21",  x"3b",  x"0b",  x"cd",  x"b9",  x"06", -- 01D8
         x"7e",  x"d3",  x"bf",  x"cd",  x"e9",  x"05",  x"cd",  x"2a", -- 01E0
         x"06",  x"23",  x"0d",  x"c2",  x"dd",  x"01",  x"cd",  x"3b", -- 01E8
         x"04",  x"11",  x"00",  x"00",  x"01",  x"3b",  x"0d",  x"c5", -- 01F0
         x"d5",  x"cd",  x"b2",  x"04",  x"d1",  x"c1",  x"7a",  x"c6", -- 01F8
         x"04",  x"fe",  x"10",  x"57",  x"c2",  x"f4",  x"01",  x"0e", -- 0200
         x"f0",  x"21",  x"10",  x"4c",  x"11",  x"20",  x"4c",  x"c5", -- 0208
         x"e5",  x"d5",  x"cd",  x"c8",  x"06",  x"cd",  x"8f",  x"05", -- 0210
         x"cd",  x"de",  x"06",  x"d1",  x"eb",  x"01",  x"20",  x"00", -- 0218
         x"09",  x"eb",  x"e1",  x"09",  x"c1",  x"0c",  x"c2",  x"0f", -- 0220
         x"02",  x"11",  x"10",  x"10",  x"01",  x"6b",  x"0d",  x"c5", -- 0228
         x"d5",  x"cd",  x"b2",  x"04",  x"d1",  x"c1",  x"7a",  x"3c", -- 0230
         x"fe",  x"20",  x"57",  x"c2",  x"2c",  x"02",  x"cd",  x"dc", -- 0238
         x"05",  x"cd",  x"2a",  x"06",  x"3e",  x"bc",  x"32",  x"8d", -- 0240
         x"e0",  x"cd",  x"04",  x"04",  x"3e",  x"bd",  x"32",  x"8d", -- 0248
         x"e0",  x"cd",  x"04",  x"04",  x"cd",  x"dc",  x"05",  x"cd", -- 0250
         x"3b",  x"04",  x"21",  x"1b",  x"0b",  x"cd",  x"1e",  x"04", -- 0258
         x"01",  x"c3",  x"08",  x"11",  x"00",  x"01",  x"cd",  x"b2", -- 0260
         x"04",  x"01",  x"f6",  x"08",  x"11",  x"00",  x"07",  x"cd", -- 0268
         x"b2",  x"04",  x"21",  x"83",  x"08",  x"1e",  x"01",  x"01", -- 0270
         x"80",  x"40",  x"cd",  x"10",  x"05",  x"cd",  x"3b",  x"04", -- 0278
         x"21",  x"af",  x"e0",  x"11",  x"bf",  x"e0",  x"0e",  x"00", -- 0280
         x"cd",  x"38",  x"08",  x"21",  x"bf",  x"e0",  x"11",  x"cf", -- 0288
         x"e0",  x"0e",  x"05",  x"cd",  x"38",  x"08",  x"21",  x"6a", -- 0290
         x"09",  x"22",  x"d0",  x"e0",  x"af",  x"32",  x"cf",  x"e0", -- 0298
         x"cd",  x"e8",  x"07",  x"cd",  x"e9",  x"05",  x"21",  x"af", -- 02A0
         x"e0",  x"11",  x"bf",  x"e0",  x"0e",  x"00",  x"cd",  x"38", -- 02A8
         x"08",  x"01",  x"da",  x"0b",  x"11",  x"00",  x"00",  x"cd", -- 02B0
         x"b2",  x"04",  x"cd",  x"12",  x"06",  x"cd",  x"26",  x"08", -- 02B8
         x"cd",  x"3b",  x"04",  x"2a",  x"d0",  x"e0",  x"7e",  x"fe", -- 02C0
         x"2e",  x"ca",  x"54",  x"03",  x"23",  x"4e",  x"eb",  x"3a", -- 02C8
         x"cf",  x"e0",  x"81",  x"fe",  x"11",  x"d2",  x"9c",  x"02", -- 02D0
         x"3a",  x"cf",  x"e0",  x"21",  x"9f",  x"e0",  x"cd",  x"b2", -- 02D8
         x"06",  x"b7",  x"3e",  x"10",  x"ca",  x"ec",  x"02",  x"2b", -- 02E0
         x"7e",  x"c6",  x"10",  x"23",  x"e5",  x"21",  x"d2",  x"e0", -- 02E8
         x"77",  x"23",  x"c6",  x"10",  x"77",  x"d6",  x"10",  x"23", -- 02F0
         x"77",  x"c6",  x"10",  x"23",  x"77",  x"e1",  x"c5",  x"d5", -- 02F8
         x"59",  x"01",  x"d2",  x"e0",  x"cd",  x"2f",  x"08",  x"d1", -- 0300
         x"c1",  x"3a",  x"cf",  x"e0",  x"21",  x"8f",  x"e0",  x"cd", -- 0308
         x"b2",  x"06",  x"b7",  x"3e",  x"10",  x"ca",  x"1d",  x"03", -- 0310
         x"2b",  x"7e",  x"c6",  x"10",  x"23",  x"e5",  x"21",  x"d2", -- 0318
         x"e0",  x"77",  x"23",  x"77",  x"c6",  x"10",  x"23",  x"77", -- 0320
         x"23",  x"77",  x"e1",  x"c5",  x"d5",  x"59",  x"01",  x"d2", -- 0328
         x"e0",  x"cd",  x"2f",  x"08",  x"d1",  x"c1",  x"21",  x"af", -- 0330
         x"e0",  x"3a",  x"cf",  x"e0",  x"cd",  x"b2",  x"06",  x"eb", -- 0338
         x"86",  x"32",  x"cf",  x"e0",  x"4e",  x"23",  x"7e",  x"12", -- 0340
         x"23",  x"13",  x"0d",  x"c2",  x"46",  x"03",  x"22",  x"d0", -- 0348
         x"e0",  x"c3",  x"c3",  x"02",  x"21",  x"8f",  x"e0",  x"01", -- 0350
         x"83",  x"08",  x"1e",  x"40",  x"cd",  x"2f",  x"08",  x"cd", -- 0358
         x"e8",  x"07",  x"21",  x"0d",  x"09",  x"cd",  x"12",  x"08", -- 0360
         x"21",  x"11",  x"09",  x"cd",  x"12",  x"08",  x"21",  x"16", -- 0368
         x"09",  x"cd",  x"12",  x"08",  x"21",  x"1d",  x"09",  x"cd", -- 0370
         x"12",  x"08",  x"06",  x"00",  x"21",  x"8f",  x"e0",  x"78", -- 0378
         x"cd",  x"b2",  x"06",  x"78",  x"2f",  x"0f",  x"0f",  x"5f", -- 0380
         x"0f",  x"57",  x"0f",  x"4f",  x"a2",  x"57",  x"79",  x"2f", -- 0388
         x"a3",  x"b2",  x"e6",  x"01",  x"ca",  x"9b",  x"03",  x"35", -- 0390
         x"c3",  x"9c",  x"03",  x"34",  x"04",  x"78",  x"fe",  x"20", -- 0398
         x"c2",  x"7c",  x"03",  x"cd",  x"e8",  x"07",  x"3a",  x"8f", -- 03A0
         x"e0",  x"fe",  x"a0",  x"c2",  x"7a",  x"03",  x"cd",  x"e9", -- 03A8
         x"05",  x"21",  x"24",  x"09",  x"cd",  x"12",  x"08",  x"cd", -- 03B0
         x"e9",  x"05",  x"21",  x"47",  x"09",  x"cd",  x"12",  x"08", -- 03B8
         x"cd",  x"e9",  x"05",  x"21",  x"af",  x"e0",  x"11",  x"bf", -- 03C0
         x"e0",  x"0e",  x"00",  x"cd",  x"38",  x"08",  x"cd",  x"e8", -- 03C8
         x"07",  x"cd",  x"3b",  x"04",  x"01",  x"01",  x"09",  x"11", -- 03D0
         x"10",  x"10",  x"cd",  x"b2",  x"04",  x"cd",  x"e9",  x"05", -- 03D8
         x"cd",  x"dc",  x"05",  x"11",  x"00",  x"00",  x"01",  x"41", -- 03E0
         x"08",  x"cd",  x"b2",  x"04",  x"14",  x"01",  x"62",  x"08", -- 03E8
         x"cd",  x"b2",  x"04",  x"14",  x"7a",  x"fe",  x"20",  x"c2", -- 03F0
         x"e6",  x"03",  x"db",  x"d1",  x"e6",  x"80",  x"c2",  x"00", -- 03F8
         x"00",  x"c3",  x"fa",  x"03",  x"0e",  x"00",  x"cd",  x"b9", -- 0400
         x"06",  x"79",  x"2f",  x"cd",  x"8c",  x"e0",  x"0c",  x"cd", -- 0408
         x"2a",  x"06",  x"c2",  x"06",  x"04",  x"cd",  x"b9",  x"06", -- 0410
         x"79",  x"2f",  x"cd",  x"8c",  x"e0",  x"c9",  x"d5",  x"c5", -- 0418
         x"01",  x"8d",  x"e0",  x"11",  x"a0",  x"10",  x"cd",  x"b9", -- 0420
         x"06",  x"7b",  x"02",  x"cd",  x"b9",  x"06",  x"7e",  x"cd", -- 0428
         x"8c",  x"e0",  x"23",  x"1c",  x"15",  x"c2",  x"29",  x"04", -- 0430
         x"c1",  x"d1",  x"c9",  x"cd",  x"c8",  x"06",  x"21",  x"00", -- 0438
         x"4c",  x"11",  x"00",  x"50",  x"0e",  x"00",  x"cd",  x"8f", -- 0440
         x"05",  x"cd",  x"de",  x"06",  x"c9",  x"06",  x"00",  x"78", -- 0448
         x"ae",  x"07",  x"47",  x"23",  x"cd",  x"5f",  x"04",  x"c2", -- 0450
         x"4f",  x"04",  x"78",  x"a9",  x"c8",  x"37",  x"c9",  x"7c", -- 0458
         x"ba",  x"c0",  x"7d",  x"bb",  x"c9",  x"4e",  x"3e",  x"01", -- 0460
         x"06",  x"08",  x"77",  x"be",  x"c4",  x"84",  x"04",  x"2f", -- 0468
         x"77",  x"be",  x"c4",  x"84",  x"04",  x"2f",  x"07",  x"05", -- 0470
         x"c2",  x"6a",  x"04",  x"71",  x"23",  x"cd",  x"5f",  x"04", -- 0478
         x"c2",  x"65",  x"04",  x"c9",  x"c5",  x"d5",  x"f5",  x"e5", -- 0480
         x"01",  x"f7",  x"0d",  x"cd",  x"ac",  x"05",  x"e1",  x"e5", -- 0488
         x"cd",  x"98",  x"04",  x"e1",  x"f1",  x"d1",  x"c1",  x"c9", -- 0490
         x"e5",  x"7c",  x"cd",  x"31",  x"05",  x"22",  x"83",  x"e0", -- 0498
         x"e1",  x"7d",  x"cd",  x"31",  x"05",  x"22",  x"85",  x"e0", -- 04A0
         x"01",  x"83",  x"e0",  x"11",  x"15",  x"10",  x"cd",  x"b2", -- 04A8
         x"04",  x"c9",  x"d5",  x"e5",  x"f5",  x"21",  x"ff",  x"4f", -- 04B0
         x"7a",  x"b7",  x"ca",  x"c9",  x"04",  x"7d",  x"d6",  x"20", -- 04B8
         x"6f",  x"7c",  x"de",  x"00",  x"67",  x"15",  x"c3",  x"b8", -- 04C0
         x"04",  x"7d",  x"93",  x"6f",  x"cd",  x"c8",  x"06",  x"cd", -- 04C8
         x"85",  x"07",  x"0a",  x"fe",  x"fe",  x"ca",  x"ea",  x"04", -- 04D0
         x"fe",  x"f2",  x"c2",  x"e4",  x"04",  x"7d",  x"f6",  x"1f", -- 04D8
         x"6f",  x"c3",  x"e5",  x"04",  x"77",  x"03",  x"23",  x"c3", -- 04E0
         x"d2",  x"04",  x"cd",  x"de",  x"06",  x"cd",  x"2a",  x"06", -- 04E8
         x"f1",  x"e1",  x"d1",  x"c9",  x"0a",  x"2f",  x"77",  x"2b", -- 04F0
         x"03",  x"1d",  x"c2",  x"f4",  x"04",  x"c9",  x"16",  x"10", -- 04F8
         x"cd",  x"85",  x"07",  x"1e",  x"40",  x"cd",  x"b9",  x"06", -- 0500
         x"cd",  x"f4",  x"04",  x"15",  x"c2",  x"03",  x"05",  x"c9", -- 0508
         x"78",  x"cd",  x"4d",  x"05",  x"32",  x"8d",  x"e0",  x"32", -- 0510
         x"8a",  x"e0",  x"cd",  x"b9",  x"06",  x"7b",  x"b7",  x"cc", -- 0518
         x"89",  x"e0",  x"7e",  x"c4",  x"8c",  x"e0",  x"cd",  x"e9", -- 0520
         x"05",  x"04",  x"78",  x"b9",  x"c8",  x"23",  x"c3",  x"10", -- 0528
         x"05",  x"d5",  x"f5",  x"e6",  x"0f",  x"21",  x"0b",  x"0b", -- 0530
         x"cd",  x"b2",  x"06",  x"56",  x"f1",  x"0f",  x"0f",  x"0f", -- 0538
         x"0f",  x"e6",  x"0f",  x"21",  x"0b",  x"0b",  x"cd",  x"b2", -- 0540
         x"06",  x"5e",  x"eb",  x"d1",  x"c9",  x"c5",  x"d5",  x"e5", -- 0548
         x"f5",  x"cd",  x"31",  x"05",  x"22",  x"80",  x"e0",  x"01", -- 0550
         x"80",  x"e0",  x"11",  x"0c",  x"07",  x"cd",  x"b2",  x"04", -- 0558
         x"f1",  x"e1",  x"d1",  x"c1",  x"c9",  x"d5",  x"e5",  x"f5", -- 0560
         x"7b",  x"3d",  x"87",  x"21",  x"87",  x"05",  x"cd",  x"b2", -- 0568
         x"06",  x"cd",  x"b9",  x"06",  x"7e",  x"d3",  x"be",  x"23", -- 0570
         x"7e",  x"d3",  x"bf",  x"21",  x"00",  x"48",  x"16",  x"20", -- 0578
         x"cd",  x"00",  x"05",  x"f1",  x"e1",  x"d1",  x"c9",  x"7d", -- 0580
         x"fe",  x"7b",  x"fb",  x"77",  x"ef",  x"6f",  x"bf",  x"cd", -- 0588
         x"85",  x"07",  x"cd",  x"8e",  x"07",  x"06",  x"40",  x"cd", -- 0590
         x"b9",  x"06",  x"79",  x"2f",  x"77",  x"2b",  x"cd",  x"5f", -- 0598
         x"04",  x"c8",  x"05",  x"c2",  x"9a",  x"05",  x"c3",  x"95", -- 05A0
         x"05",  x"01",  x"7c",  x"0d",  x"11",  x"03",  x"10",  x"cd", -- 05A8
         x"b2",  x"04",  x"cd",  x"dc",  x"05",  x"11",  x"03",  x"10", -- 05B0
         x"cd",  x"96",  x"07",  x"c9",  x"01",  x"a6",  x"0d",  x"c3", -- 05B8
         x"ac",  x"05",  x"01",  x"ba",  x"0d",  x"c3",  x"ac",  x"05", -- 05C0
         x"01",  x"93",  x"0d",  x"c3",  x"ac",  x"05",  x"f5",  x"c5", -- 05C8
         x"01",  x"4f",  x"00",  x"0b",  x"79",  x"b0",  x"c2",  x"d3", -- 05D0
         x"05",  x"c1",  x"f1",  x"c9",  x"01",  x"88",  x"13",  x"cd", -- 05D8
         x"ce",  x"05",  x"0b",  x"79",  x"b0",  x"c2",  x"df",  x"05", -- 05E0
         x"c9",  x"c5",  x"01",  x"f4",  x"01",  x"cd",  x"df",  x"05", -- 05E8
         x"c1",  x"c9",  x"32",  x"8a",  x"e0",  x"cd",  x"89",  x"e0", -- 05F0
         x"a0",  x"a9",  x"c9",  x"11",  x"88",  x"13",  x"3a",  x"88", -- 05F8
         x"e0",  x"44",  x"4d",  x"cd",  x"f2",  x"05",  x"c0",  x"cd", -- 0600
         x"ce",  x"05",  x"1b",  x"7b",  x"b2",  x"c2",  x"fe",  x"05", -- 0608
         x"37",  x"c9",  x"3e",  x"d2",  x"32",  x"88",  x"e0",  x"21", -- 0610
         x"00",  x"20",  x"cd",  x"fb",  x"05",  x"c9",  x"3e",  x"d2", -- 0618
         x"32",  x"88",  x"e0",  x"21",  x"00",  x"40",  x"cd",  x"fb", -- 0620
         x"05",  x"c9",  x"f5",  x"db",  x"d2",  x"e6",  x"40",  x"c2", -- 0628
         x"34",  x"06",  x"f1",  x"c9",  x"db",  x"d2",  x"e6",  x"40", -- 0630
         x"c2",  x"34",  x"06",  x"cd",  x"e9",  x"05",  x"db",  x"d2", -- 0638
         x"e6",  x"40",  x"ca",  x"3e",  x"06",  x"db",  x"d2",  x"e6", -- 0640
         x"40",  x"c2",  x"45",  x"06",  x"cd",  x"e9",  x"05",  x"f1", -- 0648
         x"c9",  x"3e",  x"d2",  x"32",  x"88",  x"e0",  x"21",  x"00", -- 0650
         x"10",  x"cd",  x"fb",  x"05",  x"c9",  x"cd",  x"b9",  x"06", -- 0658
         x"01",  x"05",  x"00",  x"cd",  x"df",  x"05",  x"3e",  x"d2", -- 0660
         x"01",  x"00",  x"80",  x"cd",  x"f2",  x"05",  x"37",  x"c0", -- 0668
         x"af",  x"c9",  x"e5",  x"44",  x"4d",  x"11",  x"12",  x"09", -- 0670
         x"cd",  x"b2",  x"04",  x"cd",  x"e9",  x"05",  x"01",  x"da", -- 0678
         x"0b",  x"11",  x"03",  x"0d",  x"cd",  x"b2",  x"04",  x"cd", -- 0680
         x"e9",  x"05",  x"cd",  x"12",  x"06",  x"da",  x"ac",  x"06", -- 0688
         x"16",  x"0d",  x"cd",  x"94",  x"07",  x"e1",  x"3e",  x"07", -- 0690
         x"cd",  x"b2",  x"06",  x"7e",  x"23",  x"46",  x"0e",  x"00", -- 0698
         x"cd",  x"f2",  x"05",  x"b8",  x"c8",  x"01",  x"d0",  x"0d", -- 06A0
         x"cd",  x"ac",  x"05",  x"c9",  x"cd",  x"bc",  x"05",  x"c3", -- 06A8
         x"7e",  x"06",  x"c5",  x"4f",  x"06",  x"00",  x"09",  x"c1", -- 06B0
         x"c9",  x"db",  x"d2",  x"e6",  x"80",  x"c2",  x"b9",  x"06", -- 06B8
         x"db",  x"d2",  x"e6",  x"80",  x"ca",  x"c0",  x"06",  x"c9", -- 06C0
         x"f5",  x"cd",  x"b9",  x"06",  x"3e",  x"3e",  x"d3",  x"be", -- 06C8
         x"3e",  x"ff",  x"d3",  x"bf",  x"3e",  x"04",  x"d3",  x"bd", -- 06D0
         x"3e",  x"ff",  x"d3",  x"bc",  x"f1",  x"c9",  x"f5",  x"3e", -- 06D8
         x"00",  x"d3",  x"bf",  x"3e",  x"3f",  x"d3",  x"be",  x"f1", -- 06E0
         x"c9",  x"3e",  x"38",  x"d3",  x"d7",  x"3e",  x"78",  x"d3", -- 06E8
         x"d7",  x"3e",  x"b8",  x"d3",  x"d7",  x"3e",  x"07",  x"d3", -- 06F0
         x"da",  x"3e",  x"36",  x"d3",  x"c3",  x"3e",  x"76",  x"d3", -- 06F8
         x"c3",  x"3e",  x"b8",  x"d3",  x"c3",  x"01",  x"30",  x"07", -- 0700
         x"1e",  x"09",  x"0a",  x"d5",  x"87",  x"5f",  x"16",  x"00", -- 0708
         x"21",  x"39",  x"07",  x"19",  x"5e",  x"23",  x"56",  x"7b", -- 0710
         x"d3",  x"c0",  x"7a",  x"d3",  x"c0",  x"7b",  x"d3",  x"c1", -- 0718
         x"7a",  x"d3",  x"c1",  x"d1",  x"cd",  x"e9",  x"05",  x"03", -- 0720
         x"1d",  x"cd",  x"2a",  x"06",  x"c2",  x"0a",  x"07",  x"c9", -- 0728
         x"01",  x"03",  x"05",  x"06",  x"08",  x"0a",  x"0c",  x"01", -- 0730
         x"00",  x"06",  x"00",  x"20",  x"1a",  x"a9",  x"18",  x"47", -- 0738
         x"17",  x"f8",  x"15",  x"bd",  x"14",  x"93",  x"13",  x"79", -- 0740
         x"12",  x"70",  x"11",  x"75",  x"10",  x"89",  x"0f",  x"aa", -- 0748
         x"0e",  x"d7",  x"0d",  x"21",  x"d6",  x"e0",  x"11",  x"08", -- 0750
         x"e1",  x"0e",  x"ff",  x"cd",  x"38",  x"08",  x"3e",  x"f2", -- 0758
         x"32",  x"f9",  x"e0",  x"3e",  x"fe",  x"32",  x"07",  x"e1", -- 0760
         x"32",  x"82",  x"e0",  x"32",  x"87",  x"e0",  x"3e",  x"d3", -- 0768
         x"32",  x"8c",  x"e0",  x"3e",  x"db",  x"32",  x"89",  x"e0", -- 0770
         x"3e",  x"c9",  x"32",  x"8b",  x"e0",  x"32",  x"8e",  x"e0", -- 0778
         x"3e",  x"9a",  x"d3",  x"d3",  x"c9",  x"f5",  x"7d",  x"2f", -- 0780
         x"6f",  x"7c",  x"2f",  x"67",  x"f1",  x"c9",  x"eb",  x"cd", -- 0788
         x"85",  x"07",  x"eb",  x"c9",  x"1e",  x"00",  x"01",  x"d6", -- 0790
         x"e0",  x"cd",  x"b2",  x"04",  x"c9",  x"01",  x"04",  x"00", -- 0798
         x"11",  x"00",  x"00",  x"21",  x"0b",  x"00",  x"7a",  x"c6", -- 07A0
         x"20",  x"c8",  x"57",  x"0a",  x"03",  x"c5",  x"4f",  x"cd", -- 07A8
         x"4d",  x"04",  x"c1",  x"dc",  x"b9",  x"07",  x"c3",  x"a6", -- 07B0
         x"07",  x"c5",  x"d5",  x"e5",  x"7c",  x"07",  x"07",  x"07", -- 07B8
         x"4f",  x"3a",  x"cf",  x"e0",  x"b7",  x"79",  x"ca",  x"cf", -- 07C0
         x"07",  x"32",  x"cf",  x"e0",  x"c3",  x"c9",  x"07",  x"cd", -- 07C8
         x"31",  x"05",  x"22",  x"80",  x"e0",  x"11",  x"18",  x"10", -- 07D0
         x"01",  x"80",  x"e0",  x"cd",  x"b2",  x"04",  x"01",  x"ec", -- 07D8
         x"0d",  x"cd",  x"ac",  x"05",  x"e1",  x"d1",  x"c1",  x"c9", -- 07E0
         x"c5",  x"d5",  x"e5",  x"f5",  x"cd",  x"b9",  x"06",  x"21", -- 07E8
         x"8d",  x"e0",  x"36",  x"40",  x"11",  x"8f",  x"e0",  x"0e", -- 07F0
         x"40",  x"1a",  x"2f",  x"cd",  x"8c",  x"e0",  x"13",  x"34", -- 07F8
         x"79",  x"fe",  x"20",  x"cc",  x"b9",  x"06",  x"0d",  x"c2", -- 0800
         x"f9",  x"07",  x"cd",  x"2a",  x"06",  x"f1",  x"e1",  x"d1", -- 0808
         x"c1",  x"c9",  x"4e",  x"23",  x"46",  x"23",  x"5e",  x"23", -- 0810
         x"e5",  x"c5",  x"e1",  x"c1",  x"cd",  x"2f",  x"08",  x"cd", -- 0818
         x"e8",  x"07",  x"cd",  x"e9",  x"05",  x"c9",  x"c5",  x"01", -- 0820
         x"58",  x"02",  x"cd",  x"df",  x"05",  x"c1",  x"c9",  x"0a", -- 0828
         x"77",  x"03",  x"23",  x"1d",  x"c8",  x"c3",  x"2f",  x"08", -- 0830
         x"71",  x"23",  x"cd",  x"5f",  x"04",  x"c8",  x"c3",  x"38", -- 0838
         x"08",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6", -- 0840
         x"f7",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6", -- 0848
         x"f7",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6", -- 0850
         x"f7",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6",  x"f7",  x"f6", -- 0858
         x"f7",  x"fe",  x"f8",  x"f9",  x"f8",  x"f9",  x"f8",  x"f9", -- 0860
         x"f8",  x"f9",  x"f8",  x"f9",  x"f8",  x"f9",  x"f8",  x"f9", -- 0868
         x"f8",  x"f9",  x"f8",  x"f9",  x"f8",  x"f9",  x"f8",  x"f9", -- 0870
         x"f8",  x"f9",  x"f8",  x"f9",  x"f8",  x"f9",  x"f8",  x"f9", -- 0878
         x"f8",  x"f9",  x"fe",  x"70",  x"70",  x"80",  x"80",  x"70", -- 0880
         x"70",  x"80",  x"80",  x"70",  x"70",  x"80",  x"80",  x"70", -- 0888
         x"70",  x"80",  x"80",  x"70",  x"80",  x"70",  x"80",  x"70", -- 0890
         x"80",  x"70",  x"80",  x"70",  x"80",  x"70",  x"80",  x"70", -- 0898
         x"80",  x"70",  x"80",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 08A8
         x"00",  x"00",  x"00",  x"05",  x"05",  x"05",  x"05",  x"05", -- 08B0
         x"05",  x"05",  x"05",  x"05",  x"05",  x"05",  x"05",  x"05", -- 08B8
         x"05",  x"05",  x"05",  x"a4",  x"a1",  x"9c",  x"94",  x"9e", -- 08C0
         x"a1",  x"b4",  x"a5",  x"ff",  x"a0",  x"b6",  x"b3",  x"a5", -- 08C8
         x"a3",  x"a9",  x"9c",  x"aa",  x"f2",  x"f2",  x"72",  x"9c", -- 08D0
         x"a1",  x"50",  x"b3",  x"a1",  x"9c",  x"94",  x"a5",  x"9d", -- 08D8
         x"b3",  x"9e",  x"ff",  x"a4",  x"9c",  x"a8",  x"94",  x"b3", -- 08E0
         x"95",  x"9d",  x"a6",  x"80",  x"ff",  x"9c",  x"a0",  x"89", -- 08E8
         x"9e",  x"b4",  x"a7",  x"9c",  x"94",  x"fe",  x"a7",  x"9e", -- 08F0
         x"6e",  x"a7",  x"ff",  x"a4",  x"9c",  x"a1",  x"a7",  x"a5", -- 08F8
         x"fe",  x"b4",  x"9c",  x"9d",  x"9e",  x"70",  x"ff",  x"a7", -- 0900
         x"9e",  x"6e",  x"a7",  x"a5",  x"fe",  x"af",  x"e0",  x"01", -- 0908
         x"54",  x"b3",  x"e0",  x"02",  x"65",  x"75",  x"b7",  x"e0", -- 0910
         x"04",  x"94",  x"00",  x"a4",  x"b4",  x"bb",  x"e0",  x"04", -- 0918
         x"0c",  x"1c",  x"2c",  x"5c",  x"af",  x"e0",  x"20",  x"54", -- 0920
         x"00",  x"00",  x"00",  x"75",  x"65",  x"00",  x"00",  x"00", -- 0928
         x"94",  x"b4",  x"a4",  x"1c",  x"0c",  x"5c",  x"2c",  x"09", -- 0930
         x"09",  x"09",  x"09",  x"09",  x"09",  x"09",  x"09",  x"09", -- 0938
         x"09",  x"09",  x"09",  x"09",  x"09",  x"09",  x"09",  x"af", -- 0940
         x"e0",  x"20",  x"54",  x"00",  x"00",  x"00",  x"65",  x"75", -- 0948
         x"00",  x"00",  x"a4",  x"b4",  x"94",  x"00",  x"2c",  x"5c", -- 0950
         x"0c",  x"1c",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0958
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0960
         x"07",  x"07",  x"00",  x"04",  x"00",  x"00",  x"00",  x"00", -- 0968
         x"01",  x"04",  x"00",  x"c3",  x"d3",  x"e3",  x"02",  x"04", -- 0970
         x"00",  x"a0",  x"a1",  x"a2",  x"03",  x"02",  x"4a",  x"5f", -- 0978
         x"04",  x"02",  x"4b",  x"5f",  x"05",  x"04",  x"3c",  x"4c", -- 0980
         x"4d",  x"85",  x"06",  x"01",  x"84",  x"07",  x"01",  x"f2", -- 0988
         x"08",  x"04",  x"f3",  x"80",  x"81",  x"82",  x"09",  x"04", -- 0990
         x"83",  x"90",  x"91",  x"92",  x"0a",  x"01",  x"93",  x"0b", -- 0998
         x"04",  x"a3",  x"00",  x"b3",  x"00",  x"0d",  x"01",  x"4e", -- 09A0
         x"0e",  x"01",  x"4f",  x"0f",  x"01",  x"5a",  x"10",  x"01", -- 09A8
         x"5b",  x"11",  x"01",  x"0a",  x"12",  x"01",  x"1a",  x"13", -- 09B0
         x"01",  x"2a",  x"14",  x"01",  x"3a",  x"15",  x"01",  x"0b", -- 09B8
         x"16",  x"01",  x"1b",  x"17",  x"01",  x"2b",  x"18",  x"01", -- 09C0
         x"3b",  x"19",  x"04",  x"0c",  x"1c",  x"2c",  x"5c",  x"1a", -- 09C8
         x"04",  x"0d",  x"1c",  x"1d",  x"2d",  x"1b",  x"04",  x"3d", -- 09D0
         x"1c",  x"0e",  x"1e",  x"1c",  x"04",  x"3d",  x"1c",  x"7c", -- 09D8
         x"1e",  x"1d",  x"04",  x"3e",  x"1c",  x"0f",  x"1e",  x"1e", -- 09E0
         x"04",  x"40",  x"00",  x"60",  x"70",  x"1f",  x"04",  x"41", -- 09E8
         x"51",  x"61",  x"71",  x"20",  x"04",  x"40",  x"00",  x"42", -- 09F0
         x"52",  x"21",  x"04",  x"41",  x"51",  x"62",  x"72",  x"22", -- 09F8
         x"04",  x"50",  x"53",  x"73",  x"e7",  x"23",  x"01",  x"44", -- 0A00
         x"24",  x"01",  x"54",  x"25",  x"01",  x"64",  x"26",  x"01", -- 0A08
         x"74",  x"27",  x"01",  x"45",  x"28",  x"01",  x"55",  x"29", -- 0A10
         x"01",  x"1f",  x"2a",  x"01",  x"7d",  x"2b",  x"01",  x"3f", -- 0A18
         x"2c",  x"02",  x"65",  x"75",  x"2d",  x"01",  x"46",  x"30", -- 0A20
         x"01",  x"76",  x"32",  x"04",  x"50",  x"b7",  x"73",  x"c7", -- 0A28
         x"33",  x"04",  x"56",  x"66",  x"67",  x"77",  x"34",  x"04", -- 0A30
         x"94",  x"00",  x"a4",  x"b4",  x"35",  x"04",  x"c4",  x"d4", -- 0A38
         x"e4",  x"f4",  x"36",  x"04",  x"94",  x"00",  x"95",  x"a5", -- 0A40
         x"37",  x"04",  x"c4",  x"d4",  x"86",  x"96",  x"38",  x"04", -- 0A48
         x"b5",  x"c5",  x"d5",  x"e5",  x"39",  x"04",  x"a6",  x"b6", -- 0A50
         x"c6",  x"d6",  x"3a",  x"04",  x"f5",  x"e6",  x"f6",  x"87", -- 0A58
         x"3b",  x"04",  x"00",  x"00",  x"57",  x"a7",  x"3c",  x"04", -- 0A60
         x"50",  x"b7",  x"7e",  x"7f",  x"3d",  x"01",  x"d7",  x"3e", -- 0A68
         x"02",  x"97",  x"f7",  x"3f",  x"02",  x"18",  x"28",  x"40", -- 0A70
         x"02",  x"38",  x"48",  x"41",  x"01",  x"58",  x"42",  x"01", -- 0A78
         x"68",  x"43",  x"04",  x"00",  x"00",  x"78",  x"88",  x"44", -- 0A80
         x"04",  x"00",  x"00",  x"98",  x"a8",  x"45",  x"04",  x"00", -- 0A88
         x"00",  x"b8",  x"c8",  x"46",  x"04",  x"d8",  x"00",  x"e8", -- 0A90
         x"f8",  x"47",  x"04",  x"09",  x"19",  x"29",  x"39",  x"48", -- 0A98
         x"04",  x"00",  x"49",  x"59",  x"69",  x"49",  x"04",  x"79", -- 0AA0
         x"89",  x"99",  x"a9",  x"4a",  x"04",  x"b9",  x"c9",  x"d9", -- 0AA8
         x"e9",  x"4b",  x"04",  x"5d",  x"00",  x"5e",  x"00",  x"4d", -- 0AB0
         x"01",  x"f9",  x"4e",  x"04",  x"f0",  x"1c",  x"f1",  x"2d", -- 0AB8
         x"4f",  x"02",  x"6a",  x"6b",  x"50",  x"02",  x"6c",  x"6d", -- 0AC0
         x"51",  x"04",  x"6e",  x"5d",  x"6f",  x"7a",  x"52",  x"02", -- 0AC8
         x"43",  x"63",  x"53",  x"04",  x"00",  x"00",  x"7b",  x"c8", -- 0AD0
         x"60",  x"04",  x"00",  x"47",  x"37",  x"27",  x"2e",  x"e7", -- 0AD8
         x"0a",  x"f0",  x"0a",  x"f9",  x"0a",  x"02",  x"0b",  x"94", -- 0AE0
         x"a4",  x"a1",  x"a5",  x"94",  x"9c",  x"fe",  x"d0",  x"02", -- 0AE8
         x"94",  x"96",  x"9e",  x"94",  x"9c",  x"ff",  x"fe",  x"d0", -- 0AF0
         x"20",  x"94",  x"9d",  x"b3",  x"ab",  x"ff",  x"ff",  x"fe", -- 0AF8
         x"d1",  x"20",  x"94",  x"94",  x"9e",  x"a1",  x"80",  x"ff", -- 0B00
         x"fe",  x"d1",  x"02",  x"9c",  x"a9",  x"aa",  x"ab",  x"ac", -- 0B08
         x"ad",  x"ae",  x"af",  x"b0",  x"b1",  x"a5",  x"94",  x"6e", -- 0B10
         x"f5",  x"9e",  x"f4",  x"00",  x"ef",  x"74",  x"c0",  x"d7", -- 0B18
         x"05",  x"04",  x"10",  x"23",  x"18",  x"03",  x"02",  x"28", -- 0B20
         x"24",  x"3f",  x"00",  x"01",  x"02",  x"04",  x"07",  x"08", -- 0B28
         x"10",  x"20",  x"38",  x"40",  x"80",  x"c0",  x"f8",  x"c7", -- 0B30
         x"3f",  x"00",  x"ff",  x"ff",  x"fc",  x"f3",  x"f0",  x"cf", -- 0B38
         x"cc",  x"c3",  x"c0",  x"3f",  x"3c",  x"33",  x"30",  x"0f", -- 0B40
         x"0c",  x"03",  x"00",  x"a7",  x"9e",  x"6e",  x"a7",  x"a3", -- 0B48
         x"a4",  x"a1",  x"9c",  x"9f",  x"a1",  x"a5",  x"50",  x"50", -- 0B50
         x"a5",  x"bc",  x"a4",  x"a1",  x"9c",  x"94",  x"9e",  x"a1", -- 0B58
         x"b4",  x"a5",  x"ff",  x"a0",  x"b6",  x"b3",  x"a5",  x"a3", -- 0B60
         x"a9",  x"9c",  x"9c",  x"ff",  x"f2",  x"a7",  x"9e",  x"6e", -- 0B68
         x"a7",  x"ff",  x"a4",  x"9c",  x"a1",  x"a7",  x"a5",  x"ff", -- 0B70
         x"fe",  x"a7",  x"9e",  x"6e",  x"a7",  x"ff",  x"a2",  x"ab", -- 0B78
         x"96",  x"a5",  x"ff",  x"ab",  x"94",  x"a2",  x"b4",  x"9c", -- 0B80
         x"94",  x"9c",  x"9f",  x"9c",  x"ff",  x"6e",  x"9c",  x"a4", -- 0B88
         x"a1",  x"9c",  x"94",  x"9c",  x"95",  x"a8",  x"9e",  x"a3", -- 0B90
         x"ff",  x"ff",  x"f2",  x"9d",  x"b3",  x"b8",  x"fe",  x"a7", -- 0B98
         x"9e",  x"6e",  x"a7",  x"ff",  x"a2",  x"ab",  x"96",  x"a5", -- 0BA0
         x"ff",  x"6e",  x"94",  x"b8",  x"ab",  x"b3",  x"ff",  x"6e", -- 0BA8
         x"ff",  x"a4",  x"a2",  x"96",  x"b5",  x"a7",  x"9c",  x"50", -- 0BB0
         x"fe",  x"9c",  x"a4",  x"a2",  x"6e",  x"a7",  x"b3",  x"a7", -- 0BB8
         x"9e",  x"ff",  x"50",  x"9c",  x"9d",  x"9e",  x"a7",  x"a2", -- 0BC0
         x"ff",  x"94",  x"ff",  x"50",  x"9c",  x"9d",  x"9e",  x"a7", -- 0BC8
         x"9c",  x"a4",  x"a1",  x"b3",  x"9e",  x"50",  x"9d",  x"b3", -- 0BD0
         x"b4",  x"fe",  x"9d",  x"a5",  x"95",  x"50",  x"b3",  x"a7", -- 0BD8
         x"9e",  x"ff",  x"b4",  x"9d",  x"9c",  x"a4",  x"b4",  x"a2", -- 0BE0
         x"ff",  x"a2",  x"a8",  x"a5",  x"a1",  x"fe",  x"a4",  x"a1", -- 0BE8
         x"9c",  x"94",  x"9e",  x"a1",  x"b5",  x"a7",  x"9e",  x"ff", -- 0BF0
         x"ab",  x"a5",  x"b4",  x"a1",  x"a6",  x"a7",  x"b3",  x"9e", -- 0BF8
         x"ff",  x"86",  x"9e",  x"96",  x"b3",  x"ff",  x"50",  x"9c", -- 0C00
         x"9d",  x"9e",  x"a3",  x"ff",  x"ff",  x"f2",  x"a7",  x"9c", -- 0C08
         x"a4",  x"a1",  x"b3",  x"9e",  x"50",  x"9d",  x"b3",  x"b4", -- 0C10
         x"a5",  x"fe",  x"9c",  x"a7",  x"50",  x"9e",  x"a7",  x"b5", -- 0C18
         x"a7",  x"9e",  x"ff",  x"a4",  x"9c",  x"b4",  x"a5",  x"ab", -- 0C20
         x"a5",  x"9d",  x"b3",  x"b8",  x"ff",  x"6e",  x"ac",  x"9e", -- 0C28
         x"a7",  x"ac",  x"b3",  x"b4",  x"a5",  x"ff",  x"b3",  x"9f", -- 0C30
         x"a1",  x"fe",  x"9d",  x"a5",  x"95",  x"50",  x"b3",  x"a7", -- 0C38
         x"9e",  x"ff",  x"b4",  x"9d",  x"9c",  x"a4",  x"b4",  x"a2", -- 0C40
         x"ff",  x"a0",  x"a1",  x"9c",  x"6e",  x"9c",  x"b4",  x"fe", -- 0C48
         x"ff",  x"a4",  x"a1",  x"9c",  x"94",  x"9e",  x"a1",  x"b5", -- 0C50
         x"a7",  x"9e",  x"ff",  x"a2",  x"94",  x"9e",  x"96",  x"b3", -- 0C58
         x"ac",  x"9e",  x"9d",  x"b3",  x"9e",  x"ff",  x"6e",  x"ac", -- 0C60
         x"9e",  x"a7",  x"ac",  x"b3",  x"b4",  x"a5",  x"ff",  x"ff", -- 0C68
         x"f2",  x"b3",  x"9f",  x"a1",  x"ff",  x"9d",  x"a5",  x"ff", -- 0C70
         x"a9",  x"fe",  x"a4",  x"9c",  x"94",  x"9e",  x"a1",  x"9d", -- 0C78
         x"b3",  x"a7",  x"9e",  x"ff",  x"a1",  x"a2",  x"ac",  x"b4", -- 0C80
         x"a2",  x"ff",  x"94",  x"a4",  x"a1",  x"a5",  x"94",  x"9c", -- 0C88
         x"ff",  x"a8",  x"9c",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C90
         x"ff",  x"f2",  x"ff",  x"9c",  x"a7",  x"b4",  x"a5",  x"ab", -- 0C98
         x"a5",  x"fe",  x"b4",  x"9c",  x"9d",  x"9e",  x"70",  x"ff", -- 0CA0
         x"a7",  x"9e",  x"6e",  x"a7",  x"a5",  x"ff",  x"a0",  x"b6", -- 0CA8
         x"b3",  x"a5",  x"a3",  x"a9",  x"9c",  x"9c",  x"fe",  x"a4", -- 0CB0
         x"a1",  x"9c",  x"94",  x"9e",  x"a1",  x"b4",  x"a5",  x"ff", -- 0CB8
         x"a0",  x"b6",  x"b3",  x"a5",  x"a3",  x"a9",  x"9c",  x"ab", -- 0CC0
         x"ff",  x"bc",  x"a7",  x"9e",  x"6e",  x"a7",  x"ff",  x"a4", -- 0CC8
         x"ab",  x"a2",  x"fe",  x"b4",  x"9c",  x"9d",  x"9e",  x"70", -- 0CD0
         x"ff",  x"a7",  x"9e",  x"6e",  x"a7",  x"a5",  x"ff",  x"a4", -- 0CD8
         x"ab",  x"a2",  x"bc",  x"a7",  x"9e",  x"6e",  x"a7",  x"ff", -- 0CE0
         x"9c",  x"ab",  x"a2",  x"fe",  x"b4",  x"9c",  x"9d",  x"9e", -- 0CE8
         x"70",  x"ff",  x"a7",  x"9e",  x"6e",  x"a7",  x"a5",  x"ff", -- 0CF0
         x"9c",  x"ab",  x"a2",  x"fe",  x"a4",  x"a1",  x"9c",  x"94", -- 0CF8
         x"9e",  x"a1",  x"b4",  x"a5",  x"ff",  x"a0",  x"b6",  x"b3", -- 0D00
         x"a5",  x"a3",  x"a9",  x"9c",  x"9c",  x"bb",  x"a0",  x"b6", -- 0D08
         x"b3",  x"a5",  x"a3",  x"a9",  x"9c",  x"a9",  x"ff",  x"ff", -- 0D10
         x"f2",  x"f2",  x"72",  x"9c",  x"a1",  x"50",  x"b3",  x"a1", -- 0D18
         x"9c",  x"94",  x"a5",  x"9d",  x"b3",  x"9e",  x"ff",  x"72", -- 0D20
         x"9c",  x"9d",  x"9c",  x"94",  x"a6",  x"80",  x"ff",  x"b3", -- 0D28
         x"ab",  x"9c",  x"a0",  x"a1",  x"a5",  x"95",  x"9e",  x"9d", -- 0D30
         x"b3",  x"b3",  x"fe",  x"a5",  x"a0",  x"94",  x"9f",  x"a8", -- 0D38
         x"9e",  x"95",  x"ab",  x"b3",  x"b4",  x"96",  x"50",  x"9d", -- 0D40
         x"9c",  x"a4",  x"a1",  x"6e",  x"a7",  x"a2",  x"72",  x"80", -- 0D48
         x"70",  x"ac",  x"b9",  x"86",  x"b6",  x"f2",  x"f2",  x"b7", -- 0D50
         x"b8",  x"b5",  x"89",  x"a9",  x"aa",  x"ab",  x"ac",  x"ad", -- 0D58
         x"ae",  x"af",  x"b0",  x"b1",  x"bc",  x"71",  x"a3",  x"f4", -- 0D60
         x"f5",  x"f3",  x"fe",  x"00",  x"01",  x"02",  x"03",  x"04", -- 0D68
         x"05",  x"06",  x"07",  x"08",  x"09",  x"0a",  x"0b",  x"0c", -- 0D70
         x"0d",  x"0e",  x"0f",  x"fe",  x"9c",  x"b9",  x"b3",  x"a0", -- 0D78
         x"b4",  x"a5",  x"ff",  x"50",  x"9c",  x"9d",  x"9e",  x"a7", -- 0D80
         x"9c",  x"a4",  x"a1",  x"b3",  x"9e",  x"50",  x"9d",  x"b3", -- 0D88
         x"b4",  x"a5",  x"fe",  x"9c",  x"b9",  x"b3",  x"a0",  x"b4", -- 0D90
         x"a5",  x"ff",  x"6e",  x"b3",  x"9f",  x"9d",  x"a5",  x"96", -- 0D98
         x"a5",  x"ff",  x"b4",  x"9f",  x"b3",  x"fe",  x"9c",  x"b9", -- 0DA0
         x"b3",  x"a0",  x"b4",  x"a5",  x"ff",  x"6e",  x"b3",  x"9f", -- 0DA8
         x"9d",  x"a5",  x"96",  x"a5",  x"ff",  x"a2",  x"a8",  x"a5", -- 0DB0
         x"a1",  x"fe",  x"9c",  x"b9",  x"b3",  x"a0",  x"b4",  x"a5", -- 0DB8
         x"ff",  x"6e",  x"b3",  x"9f",  x"9d",  x"a5",  x"96",  x"a5", -- 0DC0
         x"ff",  x"a0",  x"a1",  x"9c",  x"6e",  x"9c",  x"b4",  x"fe", -- 0DC8
         x"9c",  x"b9",  x"b3",  x"a0",  x"b4",  x"a5",  x"ff",  x"9d", -- 0DD0
         x"a5",  x"a4",  x"a1",  x"a5",  x"94",  x"96",  x"9e",  x"9d", -- 0DD8
         x"b3",  x"b8",  x"ff",  x"a8",  x"94",  x"b3",  x"95",  x"9e", -- 0DE0
         x"9d",  x"b3",  x"b8",  x"fe",  x"9c",  x"b9",  x"b3",  x"a0", -- 0DE8
         x"b4",  x"a5",  x"ff",  x"a4",  x"ab",  x"a2",  x"fe",  x"9c", -- 0DF0
         x"b9",  x"b3",  x"a0",  x"b4",  x"a5",  x"ff",  x"9c",  x"ab", -- 0DF8
         x"a2",  x"bc",  x"a5",  x"a8",  x"a1",  x"9e",  x"6e",  x"fe", -- 0E00
         x"cd",  x"c8",  x"06",  x"cd",  x"de",  x"06",  x"cd",  x"9d", -- 0E08
         x"07",  x"c9",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E38
         x"3e",  x"9a",  x"d3",  x"d3",  x"db",  x"d1",  x"e6",  x"80", -- 0E40
         x"c2",  x"00",  x"00",  x"31",  x"00",  x"e1",  x"01",  x"c6", -- 0E48
         x"54",  x"21",  x"76",  x"56",  x"11",  x"00",  x"f0",  x"cd", -- 0E50
         x"cd",  x"0f",  x"cd",  x"ef",  x"0f",  x"cd",  x"77",  x"14", -- 0E58
         x"cd",  x"8f",  x"14",  x"cd",  x"4f",  x"13",  x"cd",  x"6f", -- 0E60
         x"13",  x"cd",  x"f4",  x"13",  x"3e",  x"fe",  x"d3",  x"bf", -- 0E68
         x"3e",  x"7d",  x"d3",  x"be",  x"21",  x"00",  x"c0",  x"cd", -- 0E70
         x"03",  x"14",  x"cd",  x"f4",  x"13",  x"3e",  x"fb",  x"d3", -- 0E78
         x"bf",  x"3e",  x"7b",  x"d3",  x"be",  x"21",  x"00",  x"c8", -- 0E80
         x"cd",  x"03",  x"14",  x"cd",  x"f4",  x"13",  x"3e",  x"ef", -- 0E88
         x"d3",  x"bf",  x"3e",  x"77",  x"d3",  x"be",  x"21",  x"00", -- 0E90
         x"d0",  x"cd",  x"03",  x"14",  x"cd",  x"f4",  x"13",  x"3e", -- 0E98
         x"bf",  x"d3",  x"bf",  x"3e",  x"6f",  x"d3",  x"be",  x"21", -- 0EA0
         x"00",  x"d8",  x"cd",  x"03",  x"14",  x"cd",  x"6f",  x"13", -- 0EA8
         x"cd",  x"2c",  x"13",  x"cd",  x"f4",  x"13",  x"3e",  x"aa", -- 0EB0
         x"d3",  x"bf",  x"3e",  x"3f",  x"d3",  x"be",  x"af",  x"32", -- 0EB8
         x"af",  x"f0",  x"21",  x"89",  x"f0",  x"3e",  x"9c",  x"06", -- 0EC0
         x"06",  x"77",  x"23",  x"05",  x"c2",  x"c9",  x"0e",  x"01", -- 0EC8
         x"42",  x"15",  x"21",  x"47",  x"15",  x"11",  x"91",  x"f0", -- 0ED0
         x"cd",  x"cd",  x"0f",  x"11",  x"97",  x"f0",  x"cd",  x"cd", -- 0ED8
         x"0f",  x"11",  x"9d",  x"f0",  x"cd",  x"cd",  x"0f",  x"3e", -- 0EE0
         x"03",  x"32",  x"a3",  x"f0",  x"af",  x"32",  x"a4",  x"f0", -- 0EE8
         x"32",  x"a5",  x"f0",  x"3e",  x"03",  x"32",  x"a7",  x"f0", -- 0EF0
         x"3e",  x"02",  x"d3",  x"d2",  x"af",  x"32",  x"f2",  x"f0", -- 0EF8
         x"cd",  x"b3",  x"12",  x"cd",  x"7c",  x"12",  x"cd",  x"c9", -- 0F00
         x"34",  x"cd",  x"b3",  x"12",  x"cd",  x"7c",  x"12",  x"cd", -- 0F08
         x"f9",  x"34",  x"cd",  x"b3",  x"12",  x"cd",  x"7c",  x"12", -- 0F10
         x"cd",  x"2d",  x"35",  x"c3",  x"fc",  x"0e",  x"3e",  x"00", -- 0F18
         x"d3",  x"d2",  x"cd",  x"e3",  x"0f",  x"3e",  x"31",  x"32", -- 0F20
         x"a6",  x"f1",  x"3e",  x"11",  x"32",  x"ad",  x"f0",  x"cd", -- 0F28
         x"7c",  x"12",  x"cd",  x"c9",  x"34",  x"3e",  x"01",  x"32", -- 0F30
         x"ad",  x"f0",  x"cd",  x"7c",  x"12",  x"cd",  x"20",  x"37", -- 0F38
         x"3e",  x"01",  x"32",  x"af",  x"f0",  x"cd",  x"7c",  x"12", -- 0F40
         x"cd",  x"49",  x"37",  x"cd",  x"7c",  x"12",  x"cd",  x"71", -- 0F48
         x"37",  x"cd",  x"7c",  x"12",  x"cd",  x"4f",  x"38",  x"cd", -- 0F50
         x"7c",  x"12",  x"cd",  x"85",  x"45",  x"3e",  x"11",  x"32", -- 0F58
         x"ad",  x"f0",  x"cd",  x"7c",  x"12",  x"cd",  x"f9",  x"34", -- 0F60
         x"3e",  x"06",  x"32",  x"ad",  x"f0",  x"cd",  x"7c",  x"12", -- 0F68
         x"cd",  x"99",  x"38",  x"cd",  x"7c",  x"12",  x"cd",  x"b6", -- 0F70
         x"38",  x"cd",  x"7c",  x"12",  x"cd",  x"e6",  x"2c",  x"cd", -- 0F78
         x"7c",  x"12",  x"cd",  x"d3",  x"38",  x"3e",  x"11",  x"32", -- 0F80
         x"ad",  x"f0",  x"cd",  x"7c",  x"12",  x"cd",  x"c4",  x"21", -- 0F88
         x"cd",  x"bb",  x"14",  x"cd",  x"2d",  x"35",  x"3e",  x"0a", -- 0F90
         x"32",  x"ad",  x"f0",  x"cd",  x"7c",  x"12",  x"cd",  x"3d", -- 0F98
         x"2c",  x"cd",  x"7c",  x"12",  x"cd",  x"ab",  x"4b",  x"cd", -- 0FA0
         x"7c",  x"12",  x"cd",  x"3d",  x"24",  x"cd",  x"7c",  x"12", -- 0FA8
         x"cd",  x"a6",  x"4b",  x"cd",  x"7c",  x"12",  x"cd",  x"6c", -- 0FB0
         x"3f",  x"3e",  x"10",  x"32",  x"ad",  x"f0",  x"cd",  x"7c", -- 0FB8
         x"12",  x"cd",  x"46",  x"31",  x"cd",  x"7c",  x"12",  x"cd", -- 0FC0
         x"ae",  x"33",  x"c3",  x"df",  x"14",  x"c5",  x"e5",  x"0a", -- 0FC8
         x"12",  x"13",  x"78",  x"ac",  x"c2",  x"df",  x"0f",  x"79", -- 0FD0
         x"ad",  x"c2",  x"df",  x"0f",  x"e1",  x"c1",  x"c9",  x"03", -- 0FD8
         x"c3",  x"cf",  x"0f",  x"af",  x"32",  x"d6",  x"f0",  x"3c", -- 0FE0
         x"32",  x"d7",  x"f0",  x"32",  x"d9",  x"f0",  x"c9",  x"2e", -- 0FE8
         x"01",  x"26",  x"c0",  x"22",  x"d7",  x"f0",  x"24",  x"22", -- 0FF0
         x"d9",  x"f0",  x"3e",  x"38",  x"d3",  x"d7",  x"3e",  x"78", -- 0FF8
         x"d3",  x"d7",  x"3e",  x"b8",  x"d3",  x"d7",  x"3e",  x"36", -- 1000
         x"d3",  x"c3",  x"3e",  x"76",  x"d3",  x"c3",  x"3e",  x"b8", -- 1008
         x"d3",  x"c3",  x"3e",  x"07",  x"d3",  x"da",  x"af",  x"32", -- 1010
         x"d6",  x"f0",  x"c9",  x"21",  x"d7",  x"f0",  x"0e",  x"02", -- 1018
         x"35",  x"ca",  x"2b",  x"10",  x"23",  x"23",  x"0d",  x"c2", -- 1020
         x"20",  x"10",  x"c9",  x"c5",  x"e5",  x"0e",  x"0d",  x"21", -- 1028
         x"98",  x"10",  x"3a",  x"a6",  x"f1",  x"be",  x"23",  x"ca", -- 1030
         x"40",  x"10",  x"23",  x"23",  x"0d",  x"c2",  x"35",  x"10", -- 1038
         x"5e",  x"23",  x"56",  x"eb",  x"3a",  x"d6",  x"f0",  x"4f", -- 1040
         x"06",  x"00",  x"09",  x"c6",  x"02",  x"32",  x"d6",  x"f0", -- 1048
         x"7e",  x"b7",  x"ca",  x"92",  x"10",  x"57",  x"23",  x"5e", -- 1050
         x"e1",  x"72",  x"7b",  x"b7",  x"ca",  x"84",  x"10",  x"e5", -- 1058
         x"21",  x"47",  x"12",  x"16",  x"00",  x"19",  x"19",  x"5e", -- 1060
         x"23",  x"56",  x"e1",  x"23",  x"7e",  x"32",  x"01",  x"f0", -- 1068
         x"0f",  x"0f",  x"e6",  x"c0",  x"f6",  x"36",  x"d3",  x"c3", -- 1070
         x"7b",  x"cd",  x"00",  x"f0",  x"7a",  x"cd",  x"00",  x"f0", -- 1078
         x"c1",  x"c3",  x"25",  x"10",  x"23",  x"7e",  x"0f",  x"0f", -- 1080
         x"e6",  x"c0",  x"f6",  x"30",  x"d3",  x"c3",  x"c1",  x"c3", -- 1088
         x"25",  x"10",  x"32",  x"d6",  x"f0",  x"c3",  x"2d",  x"10", -- 1090
         x"47",  x"c1",  x"10",  x"4a",  x"05",  x"11",  x"42",  x"2a", -- 1098
         x"11",  x"59",  x"e2",  x"10",  x"4c",  x"f7",  x"10",  x"46", -- 10A0
         x"33",  x"11",  x"45",  x"38",  x"11",  x"57",  x"51",  x"11", -- 10A8
         x"4b",  x"5e",  x"11",  x"50",  x"a7",  x"11",  x"5a",  x"b8", -- 10B0
         x"11",  x"31",  x"f9",  x"11",  x"39",  x"1a",  x"12",  x"00", -- 10B8
         x"11",  x"03",  x"03",  x"03",  x"00",  x"04",  x"00",  x"04", -- 10C0
         x"00",  x"03",  x"0c",  x"03",  x"00",  x"04",  x"00",  x"04", -- 10C8
         x"00",  x"03",  x"08",  x"03",  x"00",  x"04",  x"00",  x"04", -- 10D0
         x"00",  x"03",  x"0c",  x"03",  x"00",  x"04",  x"00",  x"04", -- 10D8
         x"00",  x"00",  x"04",  x"01",  x"04",  x"00",  x"04",  x"05", -- 10E0
         x"04",  x"00",  x"04",  x"00",  x"04",  x"00",  x"02",  x"0d", -- 10E8
         x"02",  x"08",  x"02",  x"00",  x"02",  x"00",  x"00",  x"03", -- 10F0
         x"03",  x"03",  x"00",  x"09",  x"00",  x"09",  x"00",  x"00", -- 10F8
         x"32",  x"00",  x"32",  x"00",  x"00",  x"04",  x"01",  x"04", -- 1100
         x"00",  x"04",  x"05",  x"04",  x"00",  x"04",  x"08",  x"04", -- 1108
         x"00",  x"04",  x"0d",  x"04",  x"00",  x"04",  x"08",  x"04", -- 1110
         x"00",  x"04",  x"05",  x"04",  x"00",  x"04",  x"00",  x"04", -- 1118
         x"00",  x"06",  x"01",  x"06",  x"00",  x"04",  x"00",  x"04", -- 1120
         x"00",  x"00",  x"07",  x"05",  x"07",  x"00",  x"09",  x"01", -- 1128
         x"09",  x"00",  x"00",  x"5f",  x"0d",  x"5f",  x"00",  x"00", -- 1130
         x"06",  x"03",  x"06",  x"00",  x"06",  x"00",  x"06",  x"00", -- 1138
         x"06",  x"07",  x"06",  x"00",  x"06",  x"00",  x"06",  x"00", -- 1140
         x"06",  x"0a",  x"06",  x"0e",  x"06",  x"00",  x"06",  x"00", -- 1148
         x"00",  x"03",  x"01",  x"03",  x"00",  x"03",  x"02",  x"03", -- 1150
         x"00",  x"36",  x"00",  x"36",  x"00",  x"00",  x"06",  x"08", -- 1158
         x"06",  x"00",  x"07",  x"00",  x"07",  x"00",  x"03",  x"06", -- 1160
         x"03",  x"00",  x"03",  x"00",  x"03",  x"00",  x"03",  x"05", -- 1168
         x"03",  x"00",  x"14",  x"00",  x"14",  x"00",  x"02",  x"03", -- 1170
         x"02",  x"00",  x"06",  x"00",  x"06",  x"00",  x"02",  x"01", -- 1178
         x"02",  x"00",  x"06",  x"00",  x"06",  x"00",  x"02",  x"03", -- 1180
         x"02",  x"00",  x"06",  x"00",  x"06",  x"00",  x"02",  x"01", -- 1188
         x"02",  x"00",  x"06",  x"00",  x"06",  x"00",  x"02",  x"03", -- 1190
         x"02",  x"00",  x"06",  x"00",  x"06",  x"00",  x"02",  x"01", -- 1198
         x"02",  x"00",  x"08",  x"00",  x"08",  x"00",  x"00",  x"05", -- 11A0
         x"07",  x"05",  x"00",  x"05",  x"05",  x"05",  x"00",  x"05", -- 11A8
         x"03",  x"05",  x"00",  x"05",  x"01",  x"05",  x"00",  x"00", -- 11B0
         x"02",  x"08",  x"02",  x"00",  x"09",  x"00",  x"09",  x"00", -- 11B8
         x"04",  x"01",  x"04",  x"00",  x"07",  x"00",  x"07",  x"00", -- 11C0
         x"02",  x"01",  x"02",  x"00",  x"09",  x"00",  x"09",  x"00", -- 11C8
         x"04",  x"03",  x"04",  x"00",  x"07",  x"00",  x"07",  x"00", -- 11D0
         x"02",  x"0a",  x"02",  x"00",  x"09",  x"00",  x"09",  x"00", -- 11D8
         x"04",  x"03",  x"04",  x"00",  x"07",  x"00",  x"07",  x"00", -- 11E0
         x"02",  x"03",  x"02",  x"00",  x"09",  x"00",  x"09",  x"00", -- 11E8
         x"04",  x"01",  x"04",  x"00",  x"32",  x"00",  x"32",  x"00", -- 11F0
         x"00",  x"04",  x"04",  x"04",  x"00",  x"04",  x"09",  x"04", -- 11F8
         x"00",  x"04",  x"0b",  x"04",  x"00",  x"04",  x"09",  x"04", -- 1200
         x"00",  x"04",  x"07",  x"04",  x"00",  x"08",  x"04",  x"08", -- 1208
         x"00",  x"04",  x"10",  x"04",  x"00",  x"32",  x"00",  x"32", -- 1210
         x"00",  x"00",  x"03",  x"01",  x"03",  x"00",  x"03",  x"03", -- 1218
         x"03",  x"00",  x"03",  x"05",  x"03",  x"00",  x"03",  x"06", -- 1220
         x"03",  x"00",  x"03",  x"08",  x"03",  x"00",  x"03",  x"06", -- 1228
         x"03",  x"00",  x"03",  x"05",  x"03",  x"00",  x"03",  x"03", -- 1230
         x"03",  x"00",  x"06",  x"01",  x"06",  x"00",  x"03",  x"0d", -- 1238
         x"03",  x"00",  x"32",  x"00",  x"32",  x"00",  x"00",  x"06", -- 1240
         x"00",  x"20",  x"1a",  x"a9",  x"18",  x"47",  x"17",  x"f8", -- 1248
         x"15",  x"bd",  x"14",  x"93",  x"13",  x"79",  x"12",  x"70", -- 1250
         x"11",  x"75",  x"10",  x"89",  x"0f",  x"aa",  x"0e",  x"d7", -- 1258
         x"0d",  x"10",  x"0d",  x"50",  x"0c",  x"a4",  x"0b",  x"fc", -- 1260
         x"0a",  x"5e",  x"0a",  x"ca",  x"09",  x"57",  x"02",  x"78", -- 1268
         x"ac",  x"c2",  x"77",  x"12",  x"79",  x"ad",  x"c8",  x"03", -- 1270
         x"7a",  x"c3",  x"6e",  x"12",  x"cd",  x"77",  x"14",  x"21", -- 1278
         x"00",  x"58",  x"01",  x"00",  x"04",  x"3a",  x"ad",  x"f0", -- 1280
         x"3d",  x"ca",  x"90",  x"12",  x"09",  x"c3",  x"88",  x"12", -- 1288
         x"3a",  x"af",  x"f0",  x"b7",  x"ca",  x"9b",  x"12",  x"01", -- 1290
         x"80",  x"00",  x"09",  x"e5",  x"cd",  x"27",  x"14",  x"3a", -- 1298
         x"ad",  x"f0",  x"fe",  x"12",  x"c2",  x"ac",  x"12",  x"3e", -- 12A0
         x"01",  x"32",  x"ad",  x"f0",  x"cd",  x"fa",  x"12",  x"cd", -- 12A8
         x"8c",  x"13",  x"c9",  x"db",  x"d2",  x"e6",  x"10",  x"c2", -- 12B0
         x"f1",  x"12",  x"3e",  x"06",  x"d3",  x"c0",  x"af",  x"d3", -- 12B8
         x"c0",  x"3e",  x"06",  x"d3",  x"c1",  x"af",  x"d3",  x"c1", -- 12C0
         x"3e",  x"12",  x"32",  x"ad",  x"f0",  x"cd",  x"7c",  x"12", -- 12C8
         x"01",  x"00",  x"02",  x"db",  x"d2",  x"e6",  x"10",  x"c2", -- 12D0
         x"f1",  x"12",  x"cd",  x"8f",  x"14",  x"0b",  x"78",  x"b1", -- 12D8
         x"c2",  x"d3",  x"12",  x"3e",  x"11",  x"32",  x"ad",  x"f0", -- 12E0
         x"3e",  x"5a",  x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f", -- 12E8
         x"c9",  x"3e",  x"01",  x"32",  x"f2",  x"f0",  x"c1",  x"c3", -- 12F0
         x"1e",  x"0f",  x"3a",  x"a4",  x"f0",  x"2a",  x"8e",  x"15", -- 12F8
         x"22",  x"dd",  x"f0",  x"cd",  x"ba",  x"13",  x"3a",  x"a5", -- 1300
         x"f0",  x"2a",  x"90",  x"15",  x"22",  x"dd",  x"f0",  x"cd", -- 1308
         x"ba",  x"13",  x"3a",  x"a3",  x"f0",  x"2a",  x"92",  x"15", -- 1310
         x"22",  x"dd",  x"f0",  x"cd",  x"ba",  x"13",  x"3a",  x"ad", -- 1318
         x"f0",  x"3d",  x"2a",  x"8c",  x"15",  x"22",  x"dd",  x"f0", -- 1320
         x"cd",  x"ba",  x"13",  x"c9",  x"11",  x"7c",  x"15",  x"21", -- 1328
         x"01",  x"f0",  x"06",  x"10",  x"3e",  x"a0",  x"32",  x"01", -- 1330
         x"f0",  x"cd",  x"f4",  x"13",  x"1a",  x"cd",  x"00",  x"f0", -- 1338
         x"13",  x"34",  x"05",  x"c2",  x"3c",  x"13",  x"3e",  x"aa", -- 1340
         x"d3",  x"bf",  x"3e",  x"ff",  x"d3",  x"be",  x"c9",  x"06", -- 1348
         x"10",  x"21",  x"01",  x"f0",  x"3e",  x"a0",  x"32",  x"01", -- 1350
         x"f0",  x"cd",  x"f4",  x"13",  x"3e",  x"00",  x"cd",  x"00", -- 1358
         x"f0",  x"34",  x"05",  x"c2",  x"5e",  x"13",  x"3e",  x"aa", -- 1360
         x"d3",  x"bf",  x"3e",  x"ff",  x"d3",  x"be",  x"c9",  x"21", -- 1368
         x"00",  x"b0",  x"01",  x"00",  x"08",  x"cd",  x"9b",  x"14", -- 1370
         x"3e",  x"ff",  x"77",  x"23",  x"0b",  x"79",  x"e6",  x"1f", -- 1378
         x"c2",  x"78",  x"13",  x"cd",  x"b2",  x"14",  x"79",  x"b0", -- 1380
         x"c2",  x"75",  x"13",  x"c9",  x"3a",  x"a7",  x"f0",  x"fe", -- 1388
         x"03",  x"c8",  x"fe",  x"02",  x"ca",  x"b0",  x"13",  x"fe", -- 1390
         x"01",  x"ca",  x"a6",  x"13",  x"2a",  x"94",  x"15",  x"22", -- 1398
         x"dd",  x"f0",  x"cd",  x"e6",  x"13",  x"c9",  x"2a",  x"96", -- 13A0
         x"15",  x"22",  x"dd",  x"f0",  x"cd",  x"e6",  x"13",  x"c9", -- 13A8
         x"2a",  x"98",  x"15",  x"22",  x"dd",  x"f0",  x"cd",  x"e6", -- 13B0
         x"13",  x"c9",  x"06",  x"00",  x"32",  x"a8",  x"f0",  x"d6", -- 13B8
         x"0a",  x"da",  x"cb",  x"13",  x"04",  x"32",  x"a8",  x"f0", -- 13C0
         x"c3",  x"bf",  x"13",  x"3a",  x"a8",  x"f0",  x"5f",  x"16", -- 13C8
         x"00",  x"21",  x"24",  x"15",  x"19",  x"7e",  x"2a",  x"dd", -- 13D0
         x"f0",  x"77",  x"58",  x"21",  x"24",  x"15",  x"19",  x"7e", -- 13D8
         x"2a",  x"dd",  x"f0",  x"23",  x"77",  x"c9",  x"3e",  x"ff", -- 13E0
         x"2a",  x"dd",  x"f0",  x"06",  x"06",  x"77",  x"23",  x"05", -- 13E8
         x"c2",  x"ed",  x"13",  x"c9",  x"db",  x"d2",  x"e6",  x"80", -- 13F0
         x"c2",  x"f4",  x"13",  x"db",  x"d2",  x"e6",  x"80",  x"ca", -- 13F8
         x"fb",  x"13",  x"c9",  x"01",  x"40",  x"20",  x"11",  x"ff", -- 1400
         x"b7",  x"db",  x"d2",  x"e6",  x"80",  x"c2",  x"09",  x"14", -- 1408
         x"db",  x"d2",  x"e6",  x"80",  x"ca",  x"10",  x"14",  x"7e", -- 1410
         x"2f",  x"12",  x"1b",  x"23",  x"05",  x"c2",  x"17",  x"14", -- 1418
         x"0d",  x"c8",  x"06",  x"20",  x"c3",  x"09",  x"14",  x"3a", -- 1420
         x"af",  x"f0",  x"b7",  x"01",  x"00",  x"04",  x"1e",  x"ff", -- 1428
         x"ca",  x"38",  x"14",  x"01",  x"80",  x"03",  x"1e",  x"7f", -- 1430
         x"16",  x"b3",  x"e1",  x"e3",  x"db",  x"d2",  x"e6",  x"80", -- 1438
         x"c2",  x"3c",  x"14",  x"db",  x"d2",  x"e6",  x"80",  x"ca", -- 1440
         x"43",  x"14",  x"3e",  x"ff",  x"d3",  x"bf",  x"3e",  x"3e", -- 1448
         x"d3",  x"be",  x"7e",  x"12",  x"1b",  x"0b",  x"7d",  x"e6", -- 1450
         x"1f",  x"fe",  x"1f",  x"23",  x"ca",  x"62",  x"14",  x"c3", -- 1458
         x"52",  x"14",  x"3e",  x"aa",  x"d3",  x"bf",  x"3e",  x"3f", -- 1460
         x"d3",  x"be",  x"78",  x"b1",  x"c2",  x"3c",  x"14",  x"3a", -- 1468
         x"ad",  x"f0",  x"3c",  x"32",  x"ad",  x"f0",  x"c9",  x"cd", -- 1470
         x"f4",  x"13",  x"06",  x"10",  x"21",  x"01",  x"f0",  x"3e", -- 1478
         x"6f",  x"32",  x"01",  x"f0",  x"3e",  x"ff",  x"cd",  x"00", -- 1480
         x"f0",  x"35",  x"05",  x"c2",  x"86",  x"14",  x"c9",  x"cd", -- 1488
         x"f4",  x"13",  x"3e",  x"00",  x"d3",  x"bd",  x"3e",  x"00", -- 1490
         x"d3",  x"bc",  x"c9",  x"db",  x"d2",  x"e6",  x"80",  x"c2", -- 1498
         x"9b",  x"14",  x"db",  x"d2",  x"e6",  x"80",  x"ca",  x"a2", -- 14A0
         x"14",  x"3e",  x"ff",  x"d3",  x"bf",  x"3e",  x"3e",  x"d3", -- 14A8
         x"be",  x"c9",  x"3e",  x"aa",  x"d3",  x"bf",  x"3e",  x"3f", -- 14B0
         x"d3",  x"be",  x"c9",  x"11",  x"2e",  x"15",  x"06",  x"08", -- 14B8
         x"21",  x"09",  x"b1",  x"cd",  x"9b",  x"14",  x"1a",  x"77", -- 14C0
         x"13",  x"23",  x"05",  x"c2",  x"c6",  x"14",  x"06",  x"04", -- 14C8
         x"21",  x"14",  x"b1",  x"1a",  x"77",  x"13",  x"23",  x"05", -- 14D0
         x"c2",  x"d3",  x"14",  x"cd",  x"b2",  x"14",  x"c9",  x"11", -- 14D8
         x"36",  x"15",  x"06",  x"04",  x"21",  x"c9",  x"b1",  x"cd", -- 14E0
         x"9b",  x"14",  x"1a",  x"77",  x"13",  x"23",  x"05",  x"c2", -- 14E8
         x"ea",  x"14",  x"06",  x"08",  x"21",  x"d1",  x"b1",  x"1a", -- 14F0
         x"77",  x"13",  x"23",  x"05",  x"c2",  x"f7",  x"14",  x"cd", -- 14F8
         x"b2",  x"14",  x"3e",  x"39",  x"32",  x"a6",  x"f1",  x"af", -- 1500
         x"32",  x"f2",  x"f0",  x"3e",  x"04",  x"d3",  x"d2",  x"cd", -- 1508
         x"f4",  x"13",  x"af",  x"d3",  x"d2",  x"cd",  x"e3",  x"0f", -- 1510
         x"06",  x"ff",  x"cd",  x"9f",  x"1a",  x"05",  x"c2",  x"1a", -- 1518
         x"15",  x"c3",  x"be",  x"0e",  x"9c",  x"a9",  x"aa",  x"ab", -- 1520
         x"ac",  x"ad",  x"ae",  x"af",  x"b0",  x"b1",  x"a4",  x"a1", -- 1528
         x"b3",  x"ab",  x"9c",  x"94",  x"a5",  x"b8",  x"b3",  x"9f", -- 1530
         x"a1",  x"a5",  x"9c",  x"b4",  x"9c",  x"9d",  x"ac",  x"9e", -- 1538
         x"9d",  x"a5",  x"65",  x"64",  x"63",  x"62",  x"ff",  x"df", -- 1540
         x"fe",  x"b3",  x"fd",  x"b3",  x"e5",  x"b3",  x"e4",  x"b3", -- 1548
         x"e2",  x"b3",  x"e1",  x"b3",  x"be",  x"b3",  x"bd",  x"b3", -- 1550
         x"d2",  x"b3",  x"d1",  x"b3",  x"b2",  x"b3",  x"b1",  x"b3", -- 1558
         x"92",  x"b3",  x"91",  x"b3",  x"d0",  x"b3",  x"cf",  x"b3", -- 1560
         x"b0",  x"b3",  x"af",  x"b3",  x"90",  x"b3",  x"8f",  x"b3", -- 1568
         x"ce",  x"b3",  x"cd",  x"b3",  x"ae",  x"b3",  x"ad",  x"b3", -- 1570
         x"8e",  x"b3",  x"8d",  x"b3",  x"00",  x"ef",  x"74",  x"c0", -- 1578
         x"d7",  x"05",  x"04",  x"10",  x"23",  x"18",  x"03",  x"02", -- 1580
         x"28",  x"24",  x"3f",  x"00",  x"89",  x"f0",  x"8b",  x"f0", -- 1588
         x"8d",  x"f0",  x"8f",  x"f0",  x"91",  x"f0",  x"97",  x"f0", -- 1590
         x"9d",  x"f0",  x"46",  x"00",  x"00",  x"05",  x"57",  x"00", -- 1598
         x"00",  x"04",  x"55",  x"00",  x"00",  x"05",  x"56",  x"00", -- 15A0
         x"00",  x"30",  x"00",  x"2e",  x"01",  x"00",  x"07",  x"34", -- 15A8
         x"ff",  x"00",  x"07",  x"35",  x"08",  x"00",  x"07",  x"36", -- 15B0
         x"ff",  x"00",  x"07",  x"37",  x"08",  x"00",  x"07",  x"34", -- 15B8
         x"2f",  x"4a",  x"fe",  x"00",  x"04",  x"46",  x"f8",  x"00", -- 15C0
         x"04",  x"38",  x"fb",  x"00",  x"05",  x"39",  x"10",  x"00", -- 15C8
         x"09",  x"3a",  x"cc",  x"10",  x"f8",  x"09",  x"4d",  x"f5", -- 15D0
         x"00",  x"07",  x"38",  x"08",  x"00",  x"07",  x"46",  x"2e", -- 15D8
         x"46",  x"00",  x"00",  x"07",  x"34",  x"fd",  x"00",  x"09", -- 15E0
         x"46",  x"2e",  x"4a",  x"fe",  x"00",  x"04",  x"46",  x"fa", -- 15E8
         x"00",  x"04",  x"47",  x"04",  x"fb",  x"04",  x"47",  x"0c", -- 15F0
         x"fa",  x"04",  x"48",  x"06",  x"ff",  x"04",  x"48",  x"06", -- 15F8
         x"01",  x"04",  x"48",  x"06",  x"05",  x"04",  x"49",  x"04", -- 1600
         x"06",  x"04",  x"49",  x"0e",  x"00",  x"06",  x"4a",  x"fe", -- 1608
         x"00",  x"04",  x"46",  x"2e",  x"47",  x"0c",  x"fd",  x"08", -- 1610
         x"48",  x"05",  x"03",  x"05",  x"49",  x"00",  x"00",  x"03", -- 1618
         x"49",  x"26",  x"fe",  x"03",  x"43",  x"00",  x"02",  x"03", -- 1620
         x"44",  x"00",  x"fe",  x"03",  x"43",  x"00",  x"02",  x"03", -- 1628
         x"44",  x"00",  x"fe",  x"03",  x"43",  x"00",  x"02",  x"03", -- 1630
         x"44",  x"04",  x"09",  x"0b",  x"45",  x"00",  x"00",  x"05", -- 1638
         x"53",  x"00",  x"00",  x"05",  x"45",  x"00",  x"00",  x"05", -- 1640
         x"53",  x"00",  x"00",  x"05",  x"45",  x"00",  x"00",  x"05", -- 1648
         x"53",  x"00",  x"00",  x"05",  x"45",  x"00",  x"00",  x"05", -- 1650
         x"53",  x"00",  x"00",  x"05",  x"45",  x"00",  x"00",  x"05", -- 1658
         x"53",  x"00",  x"00",  x"05",  x"45",  x"2e",  x"4a",  x"fe", -- 1660
         x"00",  x"08",  x"46",  x"2e",  x"3c",  x"08",  x"00",  x"03", -- 1668
         x"02",  x"08",  x"00",  x"03",  x"31",  x"08",  x"00",  x"03", -- 1670
         x"01",  x"08",  x"00",  x"03",  x"3c",  x"2f",  x"fb",  x"00", -- 1678
         x"0b",  x"3b",  x"2e",  x"19",  x"00",  x"00",  x"0f",  x"1a", -- 1680
         x"00",  x"00",  x"0f",  x"4e",  x"00",  x"00",  x"0f",  x"1b", -- 1688
         x"00",  x"00",  x"0f",  x"1c",  x"00",  x"00",  x"0f",  x"1d", -- 1690
         x"00",  x"00",  x"0f",  x"1c",  x"00",  x"00",  x"0f",  x"1b", -- 1698
         x"00",  x"00",  x"0f",  x"4e",  x"00",  x"00",  x"0f",  x"1a", -- 16A0
         x"00",  x"00",  x"0f",  x"19",  x"2f",  x"25",  x"00",  x"00", -- 16A8
         x"0c",  x"26",  x"00",  x"00",  x"0c",  x"27",  x"00",  x"00", -- 16B0
         x"0c",  x"28",  x"2e",  x"49",  x"00",  x"02",  x"07",  x"44", -- 16B8
         x"cc",  x"08",  x"16",  x"07",  x"42",  x"00",  x"02",  x"01", -- 16C0
         x"43",  x"cc",  x"08",  x"16",  x"01",  x"42",  x"00",  x"04", -- 16C8
         x"01",  x"44",  x"cc",  x"08",  x"18",  x"01",  x"42",  x"2f", -- 16D0
         x"00",  x"00",  x"20",  x"00",  x"cc",  x"00",  x"00",  x"20", -- 16D8
         x"4c",  x"2e",  x"29",  x"2a",  x"2b",  x"2f",  x"00",  x"0b", -- 16E0
         x"4a",  x"fe",  x"00",  x"08",  x"46",  x"2e",  x"00",  x"00", -- 16E8
         x"09",  x"11",  x"00",  x"00",  x"09",  x"12",  x"00",  x"00", -- 16F0
         x"09",  x"13",  x"fc",  x"00",  x"09",  x"15",  x"fa",  x"00", -- 16F8
         x"09",  x"11",  x"00",  x"00",  x"09",  x"12",  x"00",  x"00", -- 1700
         x"09",  x"13",  x"00",  x"00",  x"09",  x"14",  x"fa",  x"00", -- 1708
         x"09",  x"11",  x"2f",  x"16",  x"fc",  x"00",  x"0a",  x"17", -- 1710
         x"03",  x"00",  x"06",  x"18",  x"cc",  x"f0",  x"fb",  x"06", -- 1718
         x"23",  x"2e",  x"0d",  x"fd",  x"00",  x"03",  x"0e",  x"fd", -- 1720
         x"00",  x"03",  x"0f",  x"fd",  x"ff",  x"03",  x"10",  x"fd", -- 1728
         x"00",  x"03",  x"0f",  x"fd",  x"00",  x"03",  x"0e",  x"fd", -- 1730
         x"01",  x"03",  x"0d",  x"2f",  x"06",  x"00",  x"00",  x"09", -- 1738
         x"07",  x"ff",  x"00",  x"09",  x"06",  x"fd",  x"00",  x"09", -- 1740
         x"07",  x"fc",  x"00",  x"09",  x"06",  x"fe",  x"00",  x"09", -- 1748
         x"07",  x"00",  x"00",  x"09",  x"06",  x"fe",  x"00",  x"09", -- 1750
         x"07",  x"fc",  x"00",  x"09",  x"06",  x"2f",  x"06",  x"02", -- 1758
         x"00",  x"04",  x"07",  x"02",  x"00",  x"04",  x"06",  x"02", -- 1760
         x"00",  x"04",  x"07",  x"02",  x"00",  x"04",  x"06",  x"2f", -- 1768
         x"3c",  x"00",  x"00",  x"08",  x"22",  x"00",  x"00",  x"08", -- 1770
         x"32",  x"00",  x"00",  x"08",  x"22",  x"00",  x"00",  x"08", -- 1778
         x"32",  x"00",  x"00",  x"08",  x"22",  x"00",  x"00",  x"08", -- 1780
         x"32",  x"00",  x"00",  x"08",  x"22",  x"2e",  x"01",  x"00", -- 1788
         x"00",  x"10",  x"01",  x"00",  x"00",  x"03",  x"3c",  x"00", -- 1790
         x"00",  x"03",  x"02",  x"00",  x"00",  x"03",  x"31",  x"00", -- 1798
         x"00",  x"03",  x"01",  x"00",  x"00",  x"03",  x"3c",  x"00", -- 17A0
         x"00",  x"03",  x"02",  x"00",  x"00",  x"03",  x"31",  x"00", -- 17A8
         x"00",  x"05",  x"01",  x"00",  x"00",  x"04",  x"54",  x"00", -- 17B0
         x"00",  x"04",  x"01",  x"00",  x"00",  x"04",  x"54",  x"00", -- 17B8
         x"00",  x"04",  x"01",  x"00",  x"00",  x"04",  x"54",  x"00", -- 17C0
         x"00",  x"04",  x"01",  x"00",  x"00",  x"03",  x"54",  x"00", -- 17C8
         x"00",  x"03",  x"01",  x"00",  x"00",  x"02",  x"54",  x"00", -- 17D0
         x"00",  x"02",  x"01",  x"00",  x"00",  x"02",  x"54",  x"2e", -- 17D8
         x"01",  x"01",  x"02",  x"04",  x"07",  x"03",  x"03",  x"01", -- 17E0
         x"05",  x"02",  x"07",  x"ff",  x"00",  x"04",  x"00",  x"00", -- 17E8
         x"00",  x"00",  x"01",  x"04",  x"00",  x"c3",  x"d3",  x"e3", -- 17F0
         x"02",  x"04",  x"00",  x"a0",  x"a1",  x"a2",  x"03",  x"02", -- 17F8
         x"4a",  x"5f",  x"00",  x"00",  x"04",  x"02",  x"4b",  x"5f", -- 1800
         x"00",  x"00",  x"05",  x"04",  x"3c",  x"4c",  x"4d",  x"85", -- 1808
         x"06",  x"01",  x"84",  x"00",  x"00",  x"00",  x"07",  x"01", -- 1810
         x"f2",  x"00",  x"00",  x"00",  x"08",  x"04",  x"f3",  x"80", -- 1818
         x"81",  x"82",  x"09",  x"04",  x"83",  x"90",  x"91",  x"92", -- 1820
         x"0a",  x"01",  x"93",  x"00",  x"00",  x"00",  x"0b",  x"02", -- 1828
         x"a3",  x"b3",  x"00",  x"00",  x"0d",  x"01",  x"4e",  x"00", -- 1830
         x"00",  x"00",  x"0e",  x"01",  x"4f",  x"00",  x"00",  x"00", -- 1838
         x"0f",  x"01",  x"5a",  x"00",  x"00",  x"00",  x"10",  x"01", -- 1840
         x"5b",  x"00",  x"00",  x"00",  x"11",  x"01",  x"0a",  x"00", -- 1848
         x"00",  x"00",  x"12",  x"01",  x"1a",  x"00",  x"00",  x"00", -- 1850
         x"13",  x"01",  x"2a",  x"00",  x"00",  x"00",  x"14",  x"01", -- 1858
         x"3a",  x"00",  x"00",  x"00",  x"15",  x"01",  x"0b",  x"00", -- 1860
         x"00",  x"00",  x"16",  x"01",  x"1b",  x"00",  x"00",  x"00", -- 1868
         x"17",  x"01",  x"2b",  x"00",  x"00",  x"00",  x"18",  x"01", -- 1870
         x"3b",  x"00",  x"00",  x"00",  x"19",  x"04",  x"0c",  x"1c", -- 1878
         x"2c",  x"5c",  x"1a",  x"04",  x"0d",  x"1c",  x"1d",  x"2d", -- 1880
         x"1b",  x"04",  x"3d",  x"1c",  x"0e",  x"1e",  x"1c",  x"04", -- 1888
         x"3d",  x"1c",  x"7c",  x"1e",  x"1d",  x"04",  x"3e",  x"1c", -- 1890
         x"0f",  x"1e",  x"1e",  x"04",  x"40",  x"00",  x"60",  x"70", -- 1898
         x"1f",  x"04",  x"41",  x"51",  x"61",  x"71",  x"20",  x"04", -- 18A0
         x"40",  x"00",  x"42",  x"52",  x"21",  x"04",  x"41",  x"51", -- 18A8
         x"62",  x"72",  x"22",  x"04",  x"50",  x"53",  x"73",  x"e7", -- 18B0
         x"23",  x"01",  x"44",  x"00",  x"00",  x"00",  x"24",  x"01", -- 18B8
         x"54",  x"00",  x"00",  x"00",  x"25",  x"01",  x"64",  x"00", -- 18C0
         x"00",  x"00",  x"26",  x"01",  x"74",  x"00",  x"00",  x"00", -- 18C8
         x"27",  x"01",  x"45",  x"00",  x"00",  x"00",  x"28",  x"01", -- 18D0
         x"55",  x"00",  x"00",  x"00",  x"29",  x"01",  x"1f",  x"00", -- 18D8
         x"00",  x"00",  x"2a",  x"01",  x"7d",  x"00",  x"00",  x"00", -- 18E0
         x"2b",  x"01",  x"3f",  x"00",  x"00",  x"00",  x"2c",  x"02", -- 18E8
         x"65",  x"75",  x"00",  x"00",  x"2d",  x"01",  x"46",  x"00", -- 18F0
         x"00",  x"00",  x"30",  x"01",  x"76",  x"00",  x"00",  x"00", -- 18F8
         x"31",  x"04",  x"b7",  x"50",  x"7f",  x"7e",  x"32",  x"04", -- 1900
         x"50",  x"b7",  x"73",  x"c7",  x"33",  x"04",  x"56",  x"66", -- 1908
         x"67",  x"77",  x"34",  x"04",  x"94",  x"00",  x"a4",  x"b4", -- 1910
         x"35",  x"04",  x"c4",  x"d4",  x"e4",  x"f4",  x"36",  x"04", -- 1918
         x"94",  x"00",  x"95",  x"a5",  x"37",  x"04",  x"c4",  x"d4", -- 1920
         x"86",  x"96",  x"38",  x"04",  x"b5",  x"c5",  x"d5",  x"e5", -- 1928
         x"39",  x"04",  x"a6",  x"b6",  x"c6",  x"d6",  x"3a",  x"04", -- 1930
         x"f5",  x"e6",  x"f6",  x"87",  x"3b",  x"04",  x"00",  x"00", -- 1938
         x"57",  x"a7",  x"3c",  x"04",  x"50",  x"b7",  x"7e",  x"7f", -- 1940
         x"3d",  x"01",  x"d7",  x"00",  x"00",  x"00",  x"3e",  x"03", -- 1948
         x"97",  x"f7",  x"08",  x"00",  x"3f",  x"03",  x"18",  x"28", -- 1950
         x"08",  x"00",  x"40",  x"03",  x"38",  x"48",  x"08",  x"00", -- 1958
         x"41",  x"01",  x"58",  x"00",  x"00",  x"00",  x"42",  x"01", -- 1960
         x"68",  x"00",  x"00",  x"00",  x"43",  x"04",  x"00",  x"00", -- 1968
         x"78",  x"88",  x"44",  x"04",  x"00",  x"00",  x"98",  x"a8", -- 1970
         x"45",  x"04",  x"00",  x"00",  x"b8",  x"c8",  x"46",  x"04", -- 1978
         x"d8",  x"00",  x"e8",  x"f8",  x"47",  x"04",  x"09",  x"19", -- 1980
         x"29",  x"39",  x"48",  x"04",  x"00",  x"49",  x"59",  x"69", -- 1988
         x"49",  x"04",  x"79",  x"89",  x"99",  x"a9",  x"4a",  x"04", -- 1990
         x"b9",  x"c9",  x"d9",  x"e9",  x"4b",  x"02",  x"5d",  x"5e", -- 1998
         x"00",  x"00",  x"4c",  x"01",  x"00",  x"00",  x"00",  x"00", -- 19A0
         x"4d",  x"01",  x"f9",  x"00",  x"00",  x"00",  x"4e",  x"04", -- 19A8
         x"f0",  x"1c",  x"f1",  x"2d",  x"4f",  x"02",  x"6a",  x"6b", -- 19B0
         x"00",  x"00",  x"50",  x"02",  x"6c",  x"6d",  x"00",  x"00", -- 19B8
         x"51",  x"04",  x"6e",  x"5d",  x"6f",  x"7a",  x"52",  x"02", -- 19C0
         x"43",  x"63",  x"00",  x"00",  x"53",  x"04",  x"00",  x"00", -- 19C8
         x"7b",  x"c8",  x"54",  x"04",  x"00",  x"00",  x"00",  x"93", -- 19D0
         x"55",  x"04",  x"00",  x"00",  x"79",  x"89",  x"56",  x"04", -- 19D8
         x"00",  x"00",  x"00",  x"c9",  x"57",  x"04",  x"79",  x"89", -- 19E0
         x"97",  x"f7",  x"60",  x"04",  x"00",  x"47",  x"37",  x"27", -- 19E8
         x"61",  x"03",  x"97",  x"f7",  x"58",  x"00",  x"62",  x"03", -- 19F0
         x"18",  x"28",  x"58",  x"00",  x"63",  x"03",  x"38",  x"48", -- 19F8
         x"58",  x"00",  x"64",  x"03",  x"97",  x"f7",  x"00",  x"00", -- 1A00
         x"65",  x"03",  x"18",  x"28",  x"00",  x"00",  x"66",  x"03", -- 1A08
         x"38",  x"48",  x"00",  x"00",  x"c3",  x"01",  x"b8",  x"00", -- 1A10
         x"00",  x"00",  x"c4",  x"01",  x"7b",  x"00",  x"00",  x"00", -- 1A18
         x"2f",  x"2e",  x"28",  x"37",  x"59",  x"37",  x"79",  x"37", -- 1A20
         x"57",  x"38",  x"db",  x"38",  x"a1",  x"38",  x"c6",  x"38", -- 1A28
         x"c6",  x"38",  x"4e",  x"31",  x"4e",  x"31",  x"74",  x"3f", -- 1A30
         x"b4",  x"36",  x"69",  x"3a",  x"69",  x"3a",  x"a3",  x"39", -- 1A38
         x"8c",  x"39",  x"46",  x"3a",  x"f4",  x"39",  x"f4",  x"39", -- 1A40
         x"69",  x"3a",  x"c8",  x"39",  x"46",  x"3a",  x"25",  x"42", -- 1A48
         x"eb",  x"3a",  x"eb",  x"3a",  x"a2",  x"37",  x"a3",  x"3a", -- 1A50
         x"b4",  x"3b",  x"73",  x"3b",  x"73",  x"3b",  x"64",  x"3f", -- 1A58
         x"db",  x"31",  x"41",  x"34",  x"00",  x"40",  x"21",  x"ec", -- 1A60
         x"17",  x"01",  x"05",  x"00",  x"7e",  x"fe",  x"2f",  x"c2", -- 1A68
         x"78",  x"1a",  x"31",  x"00",  x"e1",  x"c3",  x"f8",  x"0e", -- 1A70
         x"ba",  x"23",  x"ca",  x"81",  x"1a",  x"09",  x"c3",  x"6c", -- 1A78
         x"1a",  x"c9",  x"46",  x"23",  x"7e",  x"12",  x"13",  x"05", -- 1A80
         x"c2",  x"83",  x"1a",  x"c9",  x"3a",  x"a4",  x"f0",  x"e6", -- 1A88
         x"38",  x"0f",  x"0f",  x"0f",  x"47",  x"3a",  x"a4",  x"f0", -- 1A90
         x"e6",  x"0f",  x"80",  x"32",  x"05",  x"f1",  x"c9",  x"f5", -- 1A98
         x"c5",  x"d5",  x"e5",  x"3a",  x"f2",  x"f0",  x"b7",  x"ca", -- 1AA0
         x"e9",  x"1a",  x"3a",  x"a5",  x"f0",  x"fe",  x"05",  x"c2", -- 1AA8
         x"b8",  x"1a",  x"31",  x"00",  x"e1",  x"c3",  x"df",  x"14", -- 1AB0
         x"3a",  x"a6",  x"f0",  x"c6",  x"02",  x"fe",  x"64",  x"ca", -- 1AB8
         x"c8",  x"1a",  x"32",  x"a6",  x"f0",  x"c3",  x"e9",  x"1a", -- 1AC0
         x"af",  x"32",  x"a6",  x"f0",  x"3a",  x"a4",  x"f0",  x"3c", -- 1AC8
         x"32",  x"ec",  x"f0",  x"fe",  x"3c",  x"ca",  x"de",  x"1a", -- 1AD0
         x"32",  x"a4",  x"f0",  x"c3",  x"e9",  x"1a",  x"3a",  x"a5", -- 1AD8
         x"f0",  x"3c",  x"32",  x"a5",  x"f0",  x"af",  x"32",  x"a4", -- 1AE0
         x"f0",  x"3a",  x"0a",  x"f1",  x"3c",  x"32",  x"0a",  x"f1", -- 1AE8
         x"21",  x"5b",  x"f1",  x"06",  x"40",  x"11",  x"1b",  x"f1", -- 1AF0
         x"7e",  x"2f",  x"12",  x"13",  x"23",  x"05",  x"c2",  x"f8", -- 1AF8
         x"1a",  x"3a",  x"f2",  x"f0",  x"b7",  x"c2",  x"1a",  x"1b", -- 1B00
         x"db",  x"d2",  x"e6",  x"10",  x"ca",  x"1a",  x"1b",  x"31", -- 1B08
         x"00",  x"e1",  x"3e",  x"01",  x"32",  x"f2",  x"f0",  x"c3", -- 1B10
         x"1e",  x"0f",  x"db",  x"d2",  x"e6",  x"80",  x"c2",  x"1a", -- 1B18
         x"1b",  x"cd",  x"fa",  x"12",  x"cd",  x"8c",  x"13",  x"3e", -- 1B20
         x"40",  x"32",  x"4e",  x"f0",  x"cd",  x"2f",  x"f0",  x"3a", -- 1B28
         x"f2",  x"f0",  x"b7",  x"ca",  x"48",  x"1b",  x"db",  x"d1", -- 1B30
         x"e6",  x"80",  x"ca",  x"41",  x"1b",  x"31",  x"fe",  x"e0", -- 1B38
         x"c9",  x"3a",  x"a3",  x"f0",  x"b7",  x"ca",  x"b2",  x"1a", -- 1B40
         x"e1",  x"d1",  x"c1",  x"f1",  x"c9",  x"7e",  x"23",  x"c5", -- 1B48
         x"e5",  x"d5",  x"57",  x"32",  x"f9",  x"f0",  x"cd",  x"66", -- 1B50
         x"1a",  x"d1",  x"cd",  x"82",  x"1a",  x"e1",  x"c1",  x"c9", -- 1B58
         x"fe",  x"00",  x"c8",  x"0e",  x"04",  x"47",  x"1a",  x"80", -- 1B60
         x"12",  x"13",  x"0d",  x"c2",  x"66",  x"1b",  x"c9",  x"3a", -- 1B68
         x"a6",  x"f1",  x"fe",  x"45",  x"c8",  x"3a",  x"fe",  x"f0", -- 1B70
         x"b7",  x"c0",  x"3a",  x"6f",  x"f1",  x"fe",  x"d7",  x"d8", -- 1B78
         x"c1",  x"c9",  x"3a",  x"a6",  x"f1",  x"fe",  x"45",  x"c8", -- 1B80
         x"fe",  x"46",  x"ca",  x"af",  x"1d",  x"3a",  x"6f",  x"f1", -- 1B88
         x"fe",  x"f2",  x"d2",  x"a3",  x"1b",  x"fe",  x"ea",  x"da", -- 1B90
         x"9c",  x"1b",  x"c1",  x"c9",  x"fe",  x"78",  x"3e",  x"01", -- 1B98
         x"d2",  x"a4",  x"1b",  x"af",  x"32",  x"1a",  x"f1",  x"3a", -- 1BA0
         x"5f",  x"f1",  x"fe",  x"a7",  x"ca",  x"ce",  x"1b",  x"fe", -- 1BA8
         x"6f",  x"ca",  x"6c",  x"1d",  x"fe",  x"37",  x"c2",  x"d5", -- 1BB0
         x"1c",  x"3e",  x"03",  x"32",  x"e8",  x"f0",  x"3e",  x"4f", -- 1BB8
         x"32",  x"27",  x"f0",  x"32",  x"21",  x"f0",  x"3e",  x"37", -- 1BC0
         x"32",  x"24",  x"f0",  x"c3",  x"7e",  x"1d",  x"3e",  x"01", -- 1BC8
         x"32",  x"e8",  x"f0",  x"3e",  x"bf",  x"32",  x"27",  x"f0", -- 1BD0
         x"32",  x"21",  x"f0",  x"3e",  x"a7",  x"32",  x"24",  x"f0", -- 1BD8
         x"3a",  x"1a",  x"f1",  x"b7",  x"c0",  x"3a",  x"a6",  x"f1", -- 1BE0
         x"fe",  x"59",  x"ca",  x"f4",  x"1b",  x"fe",  x"42",  x"ca", -- 1BE8
         x"f4",  x"1b",  x"fe",  x"4a",  x"3a",  x"6f",  x"f1",  x"c2", -- 1BF0
         x"0d",  x"1c",  x"3a",  x"70",  x"f1",  x"fe",  x"78",  x"d2", -- 1BF8
         x"2c",  x"1d",  x"fe",  x"6d",  x"d2",  x"94",  x"1c",  x"fe", -- 1C00
         x"62",  x"d2",  x"34",  x"1c",  x"c9",  x"fe",  x"68",  x"d2", -- 1C08
         x"2c",  x"1d",  x"fe",  x"5d",  x"d2",  x"94",  x"1c",  x"fe", -- 1C10
         x"52",  x"d8",  x"3a",  x"5b",  x"f1",  x"c6",  x"18",  x"47", -- 1C18
         x"3a",  x"61",  x"f1",  x"b8",  x"c2",  x"34",  x"1c",  x"af", -- 1C20
         x"32",  x"19",  x"f1",  x"3e",  x"54",  x"32",  x"a6",  x"f1", -- 1C28
         x"cd",  x"e3",  x"0f",  x"c9",  x"00",  x"3a",  x"1a",  x"f1", -- 1C30
         x"b7",  x"3a",  x"5b",  x"f1",  x"ca",  x"42",  x"1c",  x"3a", -- 1C38
         x"5d",  x"f1",  x"cd",  x"26",  x"f0",  x"c8",  x"3a",  x"6f", -- 1C40
         x"f1",  x"fe",  x"6d",  x"da",  x"51",  x"1c",  x"fe",  x"c5", -- 1C48
         x"d8",  x"3e",  x"0a",  x"32",  x"f5",  x"f0",  x"af",  x"32", -- 1C50
         x"19",  x"f1",  x"11",  x"6f",  x"f1",  x"3a",  x"1a",  x"f1", -- 1C58
         x"b7",  x"1a",  x"ca",  x"6a",  x"1c",  x"d6",  x"d8",  x"c3", -- 1C60
         x"6c",  x"1c",  x"d6",  x"60",  x"2f",  x"3c",  x"cd",  x"60", -- 1C68
         x"1b",  x"3e",  x"02",  x"11",  x"5f",  x"f1",  x"cd",  x"60", -- 1C70
         x"1b",  x"21",  x"bb",  x"16",  x"11",  x"7f",  x"f1",  x"cd", -- 1C78
         x"4d",  x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"fa",  x"f0", -- 1C80
         x"22",  x"15",  x"f1",  x"3e",  x"46",  x"32",  x"a6",  x"f1", -- 1C88
         x"cd",  x"e3",  x"0f",  x"c9",  x"3a",  x"a6",  x"f1",  x"fe", -- 1C90
         x"54",  x"ca",  x"b8",  x"1c",  x"3a",  x"1a",  x"f1",  x"b7", -- 1C98
         x"3a",  x"5b",  x"f1",  x"ca",  x"a9",  x"1c",  x"3a",  x"5d", -- 1CA0
         x"f1",  x"cd",  x"20",  x"f0",  x"c2",  x"34",  x"1c",  x"3a", -- 1CA8
         x"5f",  x"f1",  x"cd",  x"23",  x"f0",  x"c2",  x"34",  x"1c", -- 1CB0
         x"3e",  x"01",  x"32",  x"19",  x"f1",  x"3e",  x"52",  x"32", -- 1CB8
         x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"3a",  x"0e",  x"f1", -- 1CC0
         x"32",  x"f5",  x"f0",  x"32",  x"2c",  x"f0",  x"21",  x"2a", -- 1CC8
         x"f0",  x"22",  x"15",  x"f1",  x"c9",  x"3a",  x"a6",  x"f1", -- 1CD0
         x"fe",  x"54",  x"c2",  x"f8",  x"1c",  x"af",  x"32",  x"e8", -- 1CD8
         x"f0",  x"3a",  x"1a",  x"f1",  x"b7",  x"3a",  x"6f",  x"f1", -- 1CE0
         x"c2",  x"f0",  x"1c",  x"fe",  x"5d",  x"c3",  x"f2",  x"1c", -- 1CE8
         x"fe",  x"d5",  x"d2",  x"b8",  x"1c",  x"c3",  x"fd",  x"1c", -- 1CF0
         x"fe",  x"52",  x"c2",  x"02",  x"1d",  x"af",  x"32",  x"e8", -- 1CF8
         x"f0",  x"c9",  x"fe",  x"4a",  x"c0",  x"3a",  x"e8",  x"f0", -- 1D00
         x"fe",  x"01",  x"c2",  x"1b",  x"1d",  x"3a",  x"1a",  x"f1", -- 1D08
         x"b7",  x"3a",  x"70",  x"f1",  x"c0",  x"fe",  x"78",  x"d2", -- 1D10
         x"2c",  x"1d",  x"c9",  x"fe",  x"02",  x"ca",  x"23",  x"1d", -- 1D18
         x"fe",  x"03",  x"c0",  x"3a",  x"70",  x"f1",  x"fe",  x"ef", -- 1D20
         x"d2",  x"2c",  x"1d",  x"c9",  x"af",  x"32",  x"19",  x"f1", -- 1D28
         x"32",  x"80",  x"f1",  x"32",  x"81",  x"f1",  x"32",  x"82", -- 1D30
         x"f1",  x"32",  x"8a",  x"f1",  x"3e",  x"45",  x"32",  x"a6", -- 1D38
         x"f1",  x"cd",  x"e3",  x"0f",  x"3e",  x"08",  x"11",  x"6f", -- 1D40
         x"f1",  x"cd",  x"60",  x"1b",  x"3e",  x"08",  x"11",  x"5f", -- 1D48
         x"f1",  x"cd",  x"60",  x"1b",  x"3e",  x"09",  x"32",  x"f5", -- 1D50
         x"f0",  x"21",  x"ad",  x"16",  x"11",  x"7f",  x"f1",  x"cd", -- 1D58
         x"4d",  x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"fa",  x"f0", -- 1D60
         x"22",  x"15",  x"f1",  x"c9",  x"3e",  x"02",  x"32",  x"e8", -- 1D68
         x"f0",  x"3e",  x"87",  x"32",  x"27",  x"f0",  x"32",  x"21", -- 1D70
         x"f0",  x"3e",  x"6f",  x"32",  x"24",  x"f0",  x"3a",  x"1a", -- 1D78
         x"f1",  x"b7",  x"ca",  x"34",  x"1c",  x"3a",  x"6f",  x"f1", -- 1D80
         x"fe",  x"df",  x"d2",  x"2c",  x"1d",  x"fe",  x"d5",  x"d2", -- 1D88
         x"94",  x"1c",  x"fe",  x"ca",  x"d8",  x"3a",  x"5d",  x"f1", -- 1D90
         x"c6",  x"18",  x"47",  x"3a",  x"61",  x"f1",  x"b8",  x"c2", -- 1D98
         x"34",  x"1c",  x"af",  x"32",  x"19",  x"f1",  x"3e",  x"54", -- 1DA0
         x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"c9",  x"3a", -- 1DA8
         x"5f",  x"f1",  x"fe",  x"af",  x"d8",  x"21",  x"d8",  x"16", -- 1DB0
         x"22",  x"15",  x"f1",  x"af",  x"32",  x"5f",  x"f1",  x"c9", -- 1DB8
         x"3a",  x"f4",  x"f0",  x"b7",  x"ca",  x"f1",  x"1d",  x"3a", -- 1DC0
         x"0b",  x"f1",  x"fe",  x"0c",  x"c2",  x"df",  x"1d",  x"3a", -- 1DC8
         x"78",  x"f1",  x"fe",  x"63",  x"da",  x"e7",  x"1d",  x"fe", -- 1DD0
         x"ef",  x"da",  x"f1",  x"1d",  x"c3",  x"e7",  x"1d",  x"3a", -- 1DD8
         x"78",  x"f1",  x"fe",  x"10",  x"d2",  x"f1",  x"1d",  x"af", -- 1DE0
         x"32",  x"88",  x"f1",  x"32",  x"f4",  x"f0",  x"32",  x"f3", -- 1DE8
         x"f0",  x"3a",  x"0b",  x"f1",  x"fe",  x"0c",  x"c2",  x"04", -- 1DF0
         x"1e",  x"3a",  x"e8",  x"f0",  x"fe",  x"02",  x"ca",  x"04", -- 1DF8
         x"1e",  x"fe",  x"00",  x"c0",  x"3a",  x"a6",  x"f1",  x"fe", -- 1E00
         x"45",  x"c8",  x"fe",  x"46",  x"c8",  x"fe",  x"59",  x"c2", -- 1E08
         x"17",  x"1e",  x"3a",  x"ed",  x"f0",  x"b7",  x"c0",  x"3a", -- 1E10
         x"fe",  x"f0",  x"b7",  x"ca",  x"3d",  x"1e",  x"3a",  x"ea", -- 1E18
         x"f0",  x"b7",  x"c2",  x"3d",  x"1e",  x"3a",  x"6f",  x"f1", -- 1E20
         x"47",  x"3a",  x"73",  x"f1",  x"90",  x"fa",  x"38",  x"1e", -- 1E28
         x"fe",  x"11",  x"d2",  x"3d",  x"1e",  x"c3",  x"2c",  x"1d", -- 1E30
         x"2f",  x"3c",  x"c3",  x"30",  x"1e",  x"3a",  x"a6",  x"f1", -- 1E38
         x"fe",  x"59",  x"ca",  x"ba",  x"1e",  x"3a",  x"f4",  x"f0", -- 1E40
         x"b7",  x"c8",  x"3a",  x"5f",  x"f1",  x"47",  x"3a",  x"68", -- 1E48
         x"f1",  x"90",  x"f5",  x"fe",  x"18",  x"da",  x"5a",  x"1e", -- 1E50
         x"f1",  x"c9",  x"3a",  x"fa",  x"f0",  x"fe",  x"3b",  x"c2", -- 1E58
         x"6c",  x"1e",  x"f1",  x"fe",  x"0e",  x"d8",  x"fe",  x"15", -- 1E60
         x"d0",  x"c3",  x"75",  x"1e",  x"f1",  x"f2",  x"66",  x"1e", -- 1E68
         x"2f",  x"3c",  x"fe",  x"09",  x"d0",  x"3a",  x"6f",  x"f1", -- 1E70
         x"47",  x"3a",  x"78",  x"f1",  x"90",  x"fa",  x"86",  x"1e", -- 1E78
         x"fe",  x"10",  x"d0",  x"c3",  x"2c",  x"1d",  x"2f",  x"3c", -- 1E80
         x"fe",  x"08",  x"da",  x"2c",  x"1d",  x"c9",  x"3e",  x"04", -- 1E88
         x"32",  x"f3",  x"f0",  x"32",  x"f8",  x"f0",  x"32",  x"f5", -- 1E90
         x"f0",  x"21",  x"88",  x"f1",  x"22",  x"14",  x"f0",  x"21", -- 1E98
         x"78",  x"f1",  x"22",  x"17",  x"f0",  x"21",  x"b5",  x"16", -- 1EA0
         x"11",  x"88",  x"f1",  x"cd",  x"4d",  x"1b",  x"3a",  x"f9", -- 1EA8
         x"f0",  x"32",  x"f4",  x"f0",  x"3e",  x"01",  x"32",  x"ed", -- 1EB0
         x"f0",  x"c9",  x"3a",  x"f4",  x"f0",  x"b7",  x"ca",  x"de", -- 1EB8
         x"1e",  x"3a",  x"68",  x"f1",  x"47",  x"3a",  x"6a",  x"f1", -- 1EC0
         x"b8",  x"da",  x"de",  x"1e",  x"3a",  x"7a",  x"f1",  x"47", -- 1EC8
         x"3a",  x"78",  x"f1",  x"90",  x"f2",  x"d9",  x"1e",  x"2f", -- 1ED0
         x"3c",  x"fe",  x"0f",  x"da",  x"8e",  x"1e",  x"3a",  x"fe", -- 1ED8
         x"f0",  x"b7",  x"ca",  x"45",  x"1e",  x"3a",  x"ea",  x"f0", -- 1EE0
         x"b7",  x"c2",  x"45",  x"1e",  x"3a",  x"7a",  x"f1",  x"47", -- 1EE8
         x"3a",  x"73",  x"f1",  x"90",  x"f2",  x"01",  x"1f",  x"2f", -- 1EF0
         x"3c",  x"fe",  x"18",  x"c2",  x"45",  x"1e",  x"c3",  x"06", -- 1EF8
         x"1f",  x"fe",  x"08",  x"d2",  x"45",  x"1e",  x"3e",  x"01", -- 1F00
         x"32",  x"ea",  x"f0",  x"3e",  x"08",  x"11",  x"73",  x"f1", -- 1F08
         x"cd",  x"60",  x"1b",  x"3e",  x"08",  x"11",  x"63",  x"f1", -- 1F10
         x"cd",  x"60",  x"1b",  x"3e",  x"09",  x"32",  x"f6",  x"f0", -- 1F18
         x"af",  x"32",  x"84",  x"f1",  x"32",  x"85",  x"f1",  x"32", -- 1F20
         x"86",  x"f1",  x"21",  x"ad",  x"16",  x"11",  x"83",  x"f1", -- 1F28
         x"cd",  x"4d",  x"1b",  x"3a",  x"f9",  x"f0",  x"32",  x"fe", -- 1F30
         x"f0",  x"22",  x"17",  x"f1",  x"c3",  x"45",  x"1e",  x"3a", -- 1F38
         x"87",  x"f1",  x"b7",  x"ca",  x"6a",  x"1f",  x"3a",  x"77", -- 1F40
         x"f1",  x"fe",  x"63",  x"da",  x"53",  x"1f",  x"fe",  x"e7", -- 1F48
         x"da",  x"6a",  x"1f",  x"af",  x"32",  x"87",  x"f1",  x"32", -- 1F50
         x"00",  x"f1",  x"32",  x"0a",  x"f1",  x"32",  x"eb",  x"f0", -- 1F58
         x"3c",  x"32",  x"f7",  x"f0",  x"21",  x"ee",  x"16",  x"22", -- 1F60
         x"03",  x"f1",  x"3a",  x"e8",  x"f0",  x"fe",  x"03",  x"ca", -- 1F68
         x"75",  x"1f",  x"fe",  x"00",  x"c0",  x"3a",  x"fa",  x"f0", -- 1F70
         x"fe",  x"3b",  x"3a",  x"5f",  x"f1",  x"ca",  x"86",  x"1f", -- 1F78
         x"fe",  x"3f",  x"d0",  x"c3",  x"89",  x"1f",  x"fe",  x"36", -- 1F80
         x"d0",  x"3a",  x"a6",  x"f1",  x"fe",  x"59",  x"ca",  x"af", -- 1F88
         x"1f",  x"3a",  x"00",  x"f1",  x"b7",  x"c8",  x"3a",  x"6f", -- 1F90
         x"f1",  x"47",  x"3a",  x"77",  x"f1",  x"90",  x"fa",  x"a7", -- 1F98
         x"1f",  x"fe",  x"18",  x"d0",  x"c3",  x"2c",  x"1d",  x"2f", -- 1FA0
         x"3c",  x"fe",  x"08",  x"da",  x"2c",  x"1d",  x"c9",  x"3a", -- 1FA8
         x"00",  x"f1",  x"b7",  x"ca",  x"cf",  x"1f",  x"3a",  x"ed", -- 1FB0
         x"f0",  x"b7",  x"c2",  x"cf",  x"1f",  x"3a",  x"7a",  x"f1", -- 1FB8
         x"47",  x"3a",  x"77",  x"f1",  x"90",  x"f2",  x"ca",  x"1f", -- 1FC0
         x"2f",  x"3c",  x"fe",  x"10",  x"da",  x"1d",  x"20",  x"3a", -- 1FC8
         x"ff",  x"f0",  x"b7",  x"ca",  x"91",  x"1f",  x"3a",  x"f1", -- 1FD0
         x"f0",  x"b7",  x"c2",  x"91",  x"1f",  x"3a",  x"7a",  x"f1", -- 1FD8
         x"47",  x"3a",  x"79",  x"f1",  x"90",  x"f2",  x"f2",  x"1f", -- 1FE0
         x"2f",  x"3c",  x"fe",  x"10",  x"d2",  x"91",  x"1f",  x"c3", -- 1FE8
         x"f7",  x"1f",  x"fe",  x"10",  x"d2",  x"91",  x"1f",  x"3e", -- 1FF0
         x"01",  x"32",  x"f1",  x"f0",  x"3e",  x"09",  x"32",  x"f7"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
