library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_g3 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_g3;

architecture rtl of rom_g3 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"3a",  x"a6",  x"f1",  x"fe",  x"45",  x"ca",  x"4c",  x"39", -- 0000
         x"fe",  x"46",  x"c2",  x"1b",  x"40",  x"3a",  x"5b",  x"f1", -- 0008
         x"fe",  x"c0",  x"da",  x"4c",  x"39",  x"cd",  x"2c",  x"24", -- 0010
         x"c3",  x"19",  x"3f",  x"3a",  x"1a",  x"f1",  x"b7",  x"ca", -- 0018
         x"ad",  x"40",  x"3a",  x"e8",  x"f0",  x"b7",  x"ca",  x"36", -- 0020
         x"40",  x"fe",  x"01",  x"ca",  x"6b",  x"40",  x"3a",  x"5b", -- 0028
         x"f1",  x"fe",  x"57",  x"da",  x"eb",  x"40",  x"3a",  x"6b", -- 0030
         x"f1",  x"fe",  x"27",  x"da",  x"a6",  x"3e",  x"fe",  x"34", -- 0038
         x"da",  x"53",  x"40",  x"fe",  x"38",  x"da",  x"a6",  x"3e", -- 0040
         x"fe",  x"60",  x"d2",  x"a6",  x"3e",  x"cd",  x"c4",  x"22", -- 0048
         x"c3",  x"4c",  x"39",  x"3a",  x"a6",  x"f1",  x"fe",  x"53", -- 0050
         x"ca",  x"65",  x"40",  x"fe",  x"42",  x"ca",  x"65",  x"40", -- 0058
         x"fe",  x"47",  x"c2",  x"a6",  x"3e",  x"cd",  x"a8",  x"44", -- 0060
         x"c3",  x"4c",  x"39",  x"3a",  x"6b",  x"f1",  x"fe",  x"27", -- 0068
         x"da",  x"a6",  x"3e",  x"fe",  x"34",  x"d2",  x"43",  x"40", -- 0070
         x"3a",  x"a6",  x"f1",  x"fe",  x"53",  x"ca",  x"a2",  x"40", -- 0078
         x"fe",  x"47",  x"c2",  x"a6",  x"3e",  x"3e",  x"4a",  x"32", -- 0080
         x"fa",  x"f0",  x"21",  x"66",  x"16",  x"11",  x"7b",  x"f1", -- 0088
         x"cd",  x"4d",  x"1b",  x"22",  x"15",  x"f1",  x"af",  x"32", -- 0090
         x"13",  x"f1",  x"32",  x"19",  x"f1",  x"3e",  x"01",  x"32", -- 0098
         x"f5",  x"f0",  x"3e",  x"52",  x"32",  x"a6",  x"f1",  x"cd", -- 00A0
         x"e3",  x"0f",  x"c3",  x"a6",  x"3e",  x"3a",  x"e8",  x"f0", -- 00A8
         x"b7",  x"ca",  x"c7",  x"41",  x"fe",  x"01",  x"c2",  x"c7", -- 00B0
         x"40",  x"3a",  x"6b",  x"f1",  x"fe",  x"90",  x"da",  x"4d", -- 00B8
         x"40",  x"fe",  x"e0",  x"da",  x"c7",  x"41",  x"c9",  x"3a", -- 00C0
         x"6b",  x"f1",  x"fe",  x"27",  x"da",  x"a6",  x"3e",  x"fe", -- 00C8
         x"38",  x"da",  x"65",  x"40",  x"3a",  x"9c",  x"f1",  x"b7", -- 00D0
         x"c2",  x"eb",  x"40",  x"3a",  x"6b",  x"f1",  x"fe",  x"de", -- 00D8
         x"d2",  x"4d",  x"40",  x"fe",  x"d6",  x"da",  x"a6",  x"3e", -- 00E0
         x"c3",  x"78",  x"40",  x"3a",  x"9f",  x"f1",  x"b7",  x"ca", -- 00E8
         x"76",  x"41",  x"21",  x"71",  x"f1",  x"3a",  x"6b",  x"f1", -- 00F0
         x"c6",  x"2a",  x"be",  x"da",  x"33",  x"41",  x"d6",  x"16", -- 00F8
         x"be",  x"d2",  x"33",  x"41",  x"3a",  x"61",  x"f1",  x"fe", -- 0100
         x"3e",  x"d2",  x"33",  x"41",  x"fe",  x"30",  x"da",  x"33", -- 0108
         x"41",  x"3a",  x"a6",  x"f1",  x"fe",  x"59",  x"c2",  x"33", -- 0110
         x"41",  x"3a",  x"fa",  x"f0",  x"fe",  x"39",  x"ca",  x"26", -- 0118
         x"41",  x"fe",  x"34",  x"c2",  x"33",  x"41",  x"21",  x"b6", -- 0120
         x"16",  x"22",  x"17",  x"f1",  x"af",  x"32",  x"9f",  x"f1", -- 0128
         x"c3",  x"a6",  x"3e",  x"3a",  x"6b",  x"f1",  x"d6",  x"02", -- 0130
         x"be",  x"d2",  x"76",  x"41",  x"c6",  x"18",  x"be",  x"da", -- 0138
         x"76",  x"41",  x"3a",  x"61",  x"f1",  x"fe",  x"47",  x"da", -- 0140
         x"6b",  x"41",  x"3a",  x"a6",  x"f1",  x"fe",  x"4a",  x"c2", -- 0148
         x"5f",  x"41",  x"3a",  x"fa",  x"f0",  x"fe",  x"4a",  x"ca", -- 0150
         x"5f",  x"41",  x"fe",  x"46",  x"c2",  x"76",  x"41",  x"af", -- 0158
         x"32",  x"81",  x"f1",  x"3e",  x"10",  x"32",  x"71",  x"f1", -- 0160
         x"c3",  x"4d",  x"40",  x"3a",  x"a6",  x"f1",  x"fe",  x"4c", -- 0168
         x"ca",  x"a6",  x"3e",  x"c3",  x"5f",  x"41",  x"3a",  x"6b", -- 0170
         x"f1",  x"fe",  x"ba",  x"da",  x"a6",  x"3e",  x"3a",  x"a6", -- 0178
         x"f1",  x"fe",  x"59",  x"c2",  x"bc",  x"41",  x"3a",  x"fa", -- 0180
         x"f0",  x"fe",  x"39",  x"ca",  x"93",  x"41",  x"fe",  x"3a", -- 0188
         x"c2",  x"a6",  x"3e",  x"3a",  x"74",  x"f1",  x"c6",  x"08", -- 0190
         x"32",  x"71",  x"f1",  x"3a",  x"64",  x"f1",  x"c6",  x"08", -- 0198
         x"32",  x"61",  x"f1",  x"af",  x"32",  x"9c",  x"f1",  x"32", -- 01A0
         x"81",  x"f1",  x"01",  x"84",  x"f1",  x"21",  x"87",  x"f1", -- 01A8
         x"cd",  x"6d",  x"12",  x"21",  x"b6",  x"16",  x"22",  x"17", -- 01B0
         x"f1",  x"c3",  x"4c",  x"39",  x"3a",  x"6b",  x"f1",  x"fe", -- 01B8
         x"c8",  x"da",  x"a6",  x"3e",  x"c3",  x"4d",  x"40",  x"3a", -- 01C0
         x"fa",  x"f0",  x"fe",  x"3b",  x"c2",  x"fa",  x"41",  x"21", -- 01C8
         x"6b",  x"f1",  x"3a",  x"73",  x"f1",  x"c6",  x"06",  x"be", -- 01D0
         x"da",  x"a6",  x"3e",  x"c6",  x"13",  x"be",  x"d2",  x"a6", -- 01D8
         x"3e",  x"21",  x"5d",  x"f1",  x"3a",  x"63",  x"f1",  x"d6", -- 01E0
         x"04",  x"be",  x"da",  x"a6",  x"3e",  x"c6",  x"08",  x"be", -- 01E8
         x"d2",  x"a6",  x"3e",  x"af",  x"32",  x"83",  x"f1",  x"c3", -- 01F0
         x"4d",  x"40",  x"fe",  x"46",  x"c2",  x"a6",  x"3e",  x"21", -- 01F8
         x"6b",  x"f1",  x"3a",  x"73",  x"f1",  x"c6",  x"0a",  x"be", -- 0200
         x"da",  x"a6",  x"3e",  x"c6",  x"08",  x"d2",  x"a6",  x"3e", -- 0208
         x"21",  x"5b",  x"f1",  x"3a",  x"63",  x"f1",  x"d6",  x"02", -- 0210
         x"be",  x"da",  x"a6",  x"3e",  x"d6",  x"1a",  x"be",  x"d2", -- 0218
         x"a6",  x"3e",  x"c3",  x"f3",  x"41",  x"3a",  x"1a",  x"f1", -- 0220
         x"b7",  x"ca",  x"bb",  x"42",  x"3a",  x"9e",  x"f1",  x"3d", -- 0228
         x"32",  x"9e",  x"f1",  x"cc",  x"42",  x"44",  x"3a",  x"5f", -- 0230
         x"f1",  x"fe",  x"bf",  x"c2",  x"59",  x"42",  x"3e",  x"01", -- 0238
         x"32",  x"e8",  x"f0",  x"3a",  x"a6",  x"f1",  x"fe",  x"52", -- 0240
         x"c2",  x"af",  x"42",  x"3a",  x"9d",  x"f1",  x"2f",  x"3c", -- 0248
         x"32",  x"9d",  x"f1",  x"cd",  x"47",  x"44",  x"c3",  x"bb", -- 0250
         x"42",  x"fe",  x"4f",  x"c2",  x"b7",  x"42",  x"3e",  x"03", -- 0258
         x"32",  x"e8",  x"f0",  x"3a",  x"a6",  x"f1",  x"fe",  x"52", -- 0260
         x"c2",  x"73",  x"42",  x"3e",  x"53",  x"32",  x"a6",  x"f1", -- 0268
         x"cd",  x"e3",  x"0f",  x"3a",  x"6b",  x"f1",  x"fe",  x"40", -- 0270
         x"da",  x"af",  x"42",  x"af",  x"32",  x"1a",  x"f1",  x"21", -- 0278
         x"7f",  x"8f",  x"22",  x"6f",  x"f1",  x"21",  x"87",  x"87", -- 0280
         x"22",  x"5f",  x"f1",  x"3e",  x"0a",  x"32",  x"82",  x"f1", -- 0288
         x"3e",  x"ff",  x"32",  x"9d",  x"f1",  x"21",  x"0c",  x"45", -- 0290
         x"22",  x"a7",  x"f1",  x"21",  x"e0",  x"17",  x"22",  x"06", -- 0298
         x"f1",  x"7e",  x"32",  x"e7",  x"f0",  x"af",  x"32",  x"f6", -- 02A0
         x"f0",  x"32",  x"0e",  x"f1",  x"c3",  x"bb",  x"42",  x"3e", -- 02A8
         x"08",  x"32",  x"9e",  x"f1",  x"c3",  x"bb",  x"42",  x"af", -- 02B0
         x"32",  x"e8",  x"f0",  x"3a",  x"1a",  x"f1",  x"b7",  x"c2", -- 02B8
         x"e4",  x"42",  x"3a",  x"9e",  x"f1",  x"3d",  x"32",  x"9e", -- 02C0
         x"f1",  x"cc",  x"6f",  x"44",  x"3a",  x"5f",  x"f1",  x"fe", -- 02C8
         x"bf",  x"ca",  x"d9",  x"42",  x"fe",  x"87",  x"c2",  x"e4", -- 02D0
         x"42",  x"3a",  x"9d",  x"f1",  x"2f",  x"3c",  x"32",  x"9d", -- 02D8
         x"f1",  x"cd",  x"74",  x"44",  x"3a",  x"1a",  x"f1",  x"b7", -- 02E0
         x"c2",  x"16",  x"43",  x"3a",  x"a6",  x"f1",  x"fe",  x"52", -- 02E8
         x"c2",  x"16",  x"43",  x"3a",  x"a0",  x"f1",  x"3d",  x"32", -- 02F0
         x"a0",  x"f1",  x"cc",  x"8b",  x"44",  x"af",  x"32",  x"e8", -- 02F8
         x"f0",  x"3a",  x"69",  x"f1",  x"fe",  x"bf",  x"c2",  x"16", -- 0300
         x"43",  x"3e",  x"53",  x"32",  x"a6",  x"f1",  x"cd",  x"e3", -- 0308
         x"0f",  x"3e",  x"01",  x"32",  x"e8",  x"f0",  x"3a",  x"9c", -- 0310
         x"f1",  x"b7",  x"c2",  x"33",  x"43",  x"3a",  x"9f",  x"f1", -- 0318
         x"b7",  x"ca",  x"84",  x"43",  x"3a",  x"71",  x"f1",  x"fe", -- 0320
         x"15",  x"d2",  x"33",  x"43",  x"af",  x"32",  x"9f",  x"f1", -- 0328
         x"c3",  x"84",  x"43",  x"3a",  x"a2",  x"f1",  x"b7",  x"ca", -- 0330
         x"67",  x"43",  x"3a",  x"a1",  x"f1",  x"3d",  x"32",  x"a1", -- 0338
         x"f1",  x"cc",  x"f4",  x"43",  x"3a",  x"71",  x"f1",  x"fe", -- 0340
         x"08",  x"d2",  x"84",  x"43",  x"af",  x"32",  x"a2",  x"f1", -- 0348
         x"32",  x"81",  x"f1",  x"21",  x"66",  x"56",  x"22",  x"84", -- 0350
         x"f1",  x"21",  x"77",  x"67",  x"22",  x"86",  x"f1",  x"3e", -- 0358
         x"07",  x"32",  x"a3",  x"f1",  x"c3",  x"84",  x"43",  x"3a", -- 0360
         x"a3",  x"f1",  x"3d",  x"32",  x"a3",  x"f1",  x"c2",  x"84", -- 0368
         x"43",  x"3e",  x"d7",  x"32",  x"71",  x"f1",  x"21",  x"74", -- 0370
         x"16",  x"11",  x"84",  x"f1",  x"cd",  x"4d",  x"1b",  x"3e", -- 0378
         x"01",  x"32",  x"a2",  x"f1",  x"3a",  x"1a",  x"f1",  x"b7", -- 0380
         x"c2",  x"69",  x"3a",  x"3a",  x"f6",  x"f0",  x"b7",  x"f5", -- 0388
         x"c2",  x"9d",  x"43",  x"3a",  x"0f",  x"f1",  x"3d",  x"32", -- 0390
         x"0f",  x"f1",  x"cc",  x"98",  x"23",  x"3a",  x"0e",  x"f1", -- 0398
         x"b7",  x"ca",  x"c7",  x"43",  x"f1",  x"3a",  x"73",  x"f1", -- 03A0
         x"c6",  x"03",  x"32",  x"73",  x"f1",  x"fe",  x"f3",  x"da", -- 03A8
         x"69",  x"3a",  x"af",  x"32",  x"0e",  x"f1",  x"32",  x"83", -- 03B0
         x"f1",  x"21",  x"0c",  x"45",  x"22",  x"a7",  x"f1",  x"3e", -- 03B8
         x"01",  x"32",  x"0f",  x"f1",  x"c3",  x"69",  x"3a",  x"f1", -- 03C0
         x"ca",  x"69",  x"3a",  x"3a",  x"e7",  x"f0",  x"3d",  x"32", -- 03C8
         x"e7",  x"f0",  x"c2",  x"69",  x"3a",  x"2a",  x"06",  x"f1", -- 03D0
         x"23",  x"22",  x"06",  x"f1",  x"7e",  x"fe",  x"ff",  x"ca", -- 03D8
         x"ee",  x"43",  x"c6",  x"01",  x"32",  x"e7",  x"f0",  x"af", -- 03E0
         x"32",  x"f6",  x"f0",  x"c3",  x"69",  x"3a",  x"21",  x"e0", -- 03E8
         x"17",  x"c3",  x"d9",  x"43",  x"2a",  x"17",  x"f1",  x"7e", -- 03F0
         x"fe",  x"2f",  x"ca",  x"1d",  x"44",  x"fe",  x"2e",  x"c2", -- 03F8
         x"23",  x"44",  x"3e",  x"10",  x"32",  x"9f",  x"f1",  x"32", -- 0400
         x"71",  x"f1",  x"3e",  x"4a",  x"32",  x"61",  x"f1",  x"32", -- 0408
         x"a1",  x"f1",  x"af",  x"32",  x"81",  x"f1",  x"21",  x"ca", -- 0410
         x"44",  x"22",  x"17",  x"f1",  x"c9",  x"21",  x"ca",  x"44", -- 0418
         x"22",  x"17",  x"f1",  x"3a",  x"71",  x"f1",  x"86",  x"32", -- 0420
         x"71",  x"f1",  x"23",  x"3a",  x"61",  x"f1",  x"86",  x"32", -- 0428
         x"61",  x"f1",  x"23",  x"7e",  x"32",  x"a1",  x"f1",  x"23", -- 0430
         x"11",  x"81",  x"f1",  x"cd",  x"4d",  x"1b",  x"22",  x"17", -- 0438
         x"f1",  x"c9",  x"3e",  x"01",  x"32",  x"9e",  x"f1",  x"3a", -- 0440
         x"a6",  x"f1",  x"fe",  x"52",  x"c2",  x"67",  x"44",  x"21", -- 0448
         x"6a",  x"f1",  x"3a",  x"9d",  x"f1",  x"86",  x"77",  x"06", -- 0450
         x"06",  x"21",  x"5b",  x"f1",  x"3a",  x"9d",  x"f1",  x"86", -- 0458
         x"77",  x"23",  x"05",  x"c2",  x"5c",  x"44",  x"c9",  x"06", -- 0460
         x"02",  x"21",  x"5f",  x"f1",  x"c3",  x"5c",  x"44",  x"3e", -- 0468
         x"01",  x"32",  x"9e",  x"f1",  x"06",  x"03",  x"21",  x"5f", -- 0470
         x"f1",  x"3a",  x"9d",  x"f1",  x"86",  x"77",  x"23",  x"05", -- 0478
         x"c8",  x"78",  x"fe",  x"01",  x"c2",  x"79",  x"44",  x"23", -- 0480
         x"c3",  x"79",  x"44",  x"3e",  x"01",  x"32",  x"a0",  x"f1", -- 0488
         x"01",  x"02",  x"04",  x"11",  x"5b",  x"f1",  x"1a",  x"3c", -- 0490
         x"12",  x"13",  x"05",  x"c2",  x"96",  x"44",  x"0d",  x"c8", -- 0498
         x"06",  x"03",  x"11",  x"68",  x"f1",  x"c3",  x"96",  x"44", -- 04A0
         x"af",  x"32",  x"13",  x"f1",  x"32",  x"14",  x"f1",  x"3e", -- 04A8
         x"46",  x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"21", -- 04B0
         x"c4",  x"44",  x"22",  x"15",  x"f1",  x"3e",  x"01",  x"32", -- 04B8
         x"f5",  x"f0",  x"c9",  x"46",  x"00",  x"06",  x"05",  x"46", -- 04C0
         x"2f",  x"29",  x"fa",  x"ff",  x"09",  x"2a",  x"fa",  x"fd", -- 04C8
         x"09",  x"2b",  x"fa",  x"fa",  x"09",  x"29",  x"fa",  x"fa", -- 04D0
         x"09",  x"2a",  x"fa",  x"fa",  x"09",  x"2b",  x"fa",  x"fa", -- 04D8
         x"09",  x"29",  x"fa",  x"fd",  x"09",  x"2a",  x"fa",  x"ff", -- 04E0
         x"09",  x"2b",  x"fa",  x"01",  x"09",  x"29",  x"fa",  x"03", -- 04E8
         x"09",  x"2a",  x"fa",  x"06",  x"09",  x"2b",  x"fa",  x"06", -- 04F0
         x"09",  x"29",  x"fa",  x"06",  x"09",  x"2a",  x"fa",  x"06", -- 04F8
         x"09",  x"2b",  x"fa",  x"03",  x"09",  x"29",  x"fa",  x"01", -- 0500
         x"09",  x"2b",  x"2f",  x"11",  x"fc",  x"00",  x"09",  x"16", -- 0508
         x"04",  x"00",  x"0a",  x"17",  x"cc",  x"fd",  x"00",  x"09", -- 0510
         x"18",  x"03",  x"00",  x"04",  x"11",  x"2e",  x"3a",  x"19", -- 0518
         x"f1",  x"b7",  x"ca",  x"4c",  x"39",  x"79",  x"fe",  x"4c", -- 0520
         x"c2",  x"35",  x"45",  x"af",  x"32",  x"13",  x"f1",  x"32", -- 0528
         x"19",  x"f1",  x"c3",  x"10",  x"3e",  x"fe",  x"53",  x"c2", -- 0530
         x"62",  x"45",  x"3a",  x"fa",  x"f0",  x"fe",  x"46",  x"ca", -- 0538
         x"4c",  x"39",  x"21",  x"66",  x"16",  x"11",  x"7b",  x"f1", -- 0540
         x"cd",  x"4d",  x"1b",  x"22",  x"15",  x"f1",  x"3e",  x"02", -- 0548
         x"32",  x"f5",  x"f0",  x"3e",  x"4a",  x"32",  x"fa",  x"f0", -- 0550
         x"af",  x"32",  x"13",  x"f1",  x"32",  x"19",  x"f1",  x"c3", -- 0558
         x"4c",  x"39",  x"fe",  x"59",  x"c2",  x"4c",  x"39",  x"3a", -- 0560
         x"fa",  x"f0",  x"fe",  x"46",  x"c2",  x"7f",  x"45",  x"21", -- 0568
         x"c6",  x"15",  x"22",  x"15",  x"f1",  x"af",  x"32",  x"13", -- 0570
         x"f1",  x"32",  x"19",  x"f1",  x"c3",  x"5d",  x"3c",  x"21", -- 0578
         x"c1",  x"15",  x"c3",  x"45",  x"45",  x"21",  x"d0",  x"49", -- 0580
         x"3e",  x"05",  x"32",  x"0b",  x"f1",  x"3e",  x"01",  x"32", -- 0588
         x"ec",  x"f0",  x"cd",  x"7c",  x"49",  x"21",  x"63",  x"4b", -- 0590
         x"cd",  x"7c",  x"49",  x"cd",  x"9f",  x"1a",  x"21",  x"c8", -- 0598
         x"f0",  x"3e",  x"08",  x"cd",  x"62",  x"48",  x"21",  x"b4", -- 05A0
         x"f0",  x"af",  x"cd",  x"62",  x"48",  x"cd",  x"9f",  x"1a", -- 05A8
         x"d2",  x"9e",  x"45",  x"af",  x"32",  x"19",  x"f1",  x"32", -- 05B0
         x"b3",  x"f0",  x"3e",  x"ff",  x"32",  x"b0",  x"f0",  x"3e", -- 05B8
         x"53",  x"32",  x"a6",  x"f1",  x"af",  x"32",  x"b1",  x"f0", -- 05C0
         x"cd",  x"9f",  x"1a",  x"3a",  x"b3",  x"f0",  x"b7",  x"c2", -- 05C8
         x"d9",  x"45",  x"21",  x"c0",  x"f0",  x"af",  x"cd",  x"62", -- 05D0
         x"48",  x"3a",  x"a6",  x"f1",  x"fe",  x"59",  x"c2",  x"10", -- 05D8
         x"46",  x"3a",  x"ba",  x"f0",  x"fe",  x"14",  x"c2",  x"10", -- 05E0
         x"46",  x"21",  x"c4",  x"f0",  x"3e",  x"0a",  x"cd",  x"62", -- 05E8
         x"48",  x"cd",  x"9f",  x"1a",  x"d2",  x"e9",  x"45",  x"3a", -- 05F0
         x"6b",  x"f1",  x"4f",  x"3a",  x"75",  x"f1",  x"c6",  x"0a", -- 05F8
         x"cd",  x"93",  x"49",  x"fe",  x"0b",  x"da",  x"dc",  x"47", -- 0600
         x"3e",  x"04",  x"32",  x"95",  x"f1",  x"c3",  x"a1",  x"46", -- 0608
         x"3a",  x"b1",  x"f0",  x"b7",  x"ca",  x"2d",  x"46",  x"3a", -- 0610
         x"6f",  x"f1",  x"32",  x"73",  x"f1",  x"c6",  x"10",  x"32", -- 0618
         x"74",  x"f1",  x"3a",  x"5f",  x"f1",  x"c6",  x"05",  x"32", -- 0620
         x"63",  x"f1",  x"32",  x"64",  x"f1",  x"21",  x"c8",  x"f0", -- 0628
         x"3e",  x"08",  x"cd",  x"62",  x"48",  x"3a",  x"b0",  x"f0", -- 0630
         x"b7",  x"ca",  x"51",  x"46",  x"21",  x"b8",  x"f0",  x"3e", -- 0638
         x"04",  x"cd",  x"62",  x"48",  x"d2",  x"51",  x"46",  x"af", -- 0640
         x"32",  x"b0",  x"f0",  x"32",  x"19",  x"f1",  x"32",  x"a6", -- 0648
         x"f1",  x"3a",  x"5f",  x"f1",  x"6f",  x"3a",  x"6b",  x"f1", -- 0650
         x"4f",  x"3a",  x"6f",  x"f1",  x"fe",  x"e8",  x"d2",  x"96", -- 0658
         x"46",  x"c6",  x"0a",  x"67",  x"cd",  x"93",  x"49",  x"fe", -- 0660
         x"05",  x"da",  x"05",  x"47",  x"3a",  x"73",  x"f1",  x"c6", -- 0668
         x"08",  x"4c",  x"cd",  x"93",  x"49",  x"fe",  x"07",  x"d2", -- 0670
         x"7d",  x"46",  x"c3",  x"8e",  x"46",  x"3a",  x"19",  x"f1", -- 0678
         x"b7",  x"c2",  x"c8",  x"45",  x"cd",  x"b6",  x"20",  x"cd", -- 0680
         x"98",  x"49",  x"da",  x"c8",  x"45",  x"e9",  x"3e",  x"ff", -- 0688
         x"32",  x"b1",  x"f0",  x"c3",  x"7d",  x"46",  x"3a",  x"b1", -- 0690
         x"f0",  x"b7",  x"c0",  x"3a",  x"6f",  x"f1",  x"c3",  x"61", -- 0698
         x"46",  x"cd",  x"1a",  x"48",  x"3e",  x"53",  x"32",  x"a6", -- 06A0
         x"f1",  x"21",  x"6d",  x"4a",  x"22",  x"b8",  x"f0",  x"21", -- 06A8
         x"00",  x"00",  x"22",  x"ba",  x"f0",  x"c3",  x"c8",  x"45", -- 06B0
         x"3a",  x"a6",  x"f1",  x"fe",  x"47",  x"ca",  x"c8",  x"45", -- 06B8
         x"cd",  x"1a",  x"48",  x"3e",  x"47",  x"32",  x"a6",  x"f1", -- 06C0
         x"21",  x"73",  x"4a",  x"c3",  x"ac",  x"46",  x"3a",  x"a6", -- 06C8
         x"f1",  x"fe",  x"42",  x"ca",  x"c8",  x"45",  x"cd",  x"1a", -- 06D0
         x"48",  x"3e",  x"42",  x"32",  x"a6",  x"f1",  x"21",  x"85", -- 06D8
         x"4a",  x"c3",  x"ac",  x"46",  x"cd",  x"1a",  x"48",  x"3e", -- 06E0
         x"4c",  x"32",  x"a6",  x"f1",  x"21",  x"8f",  x"4a",  x"c3", -- 06E8
         x"ac",  x"46",  x"3e",  x"ff",  x"32",  x"b0",  x"f0",  x"32", -- 06F0
         x"19",  x"f1",  x"3e",  x"4a",  x"32",  x"a6",  x"f1",  x"21", -- 06F8
         x"95",  x"4a",  x"c3",  x"ac",  x"46",  x"3a",  x"b3",  x"f0", -- 0700
         x"b7",  x"c2",  x"7d",  x"46",  x"01",  x"7b",  x"f1",  x"1e", -- 0708
         x"08",  x"cd",  x"ef",  x"48",  x"2a",  x"6b",  x"f1",  x"22", -- 0710
         x"76",  x"f1",  x"2a",  x"6d",  x"f1",  x"22",  x"78",  x"f1", -- 0718
         x"2a",  x"5b",  x"f1",  x"22",  x"66",  x"f1",  x"2a",  x"5d", -- 0720
         x"f1",  x"22",  x"68",  x"f1",  x"3a",  x"76",  x"f1",  x"d6", -- 0728
         x"19",  x"32",  x"75",  x"f1",  x"3a",  x"66",  x"f1",  x"c6", -- 0730
         x"10",  x"32",  x"65",  x"f1",  x"3e",  x"68",  x"32",  x"85", -- 0738
         x"f1",  x"3e",  x"05",  x"32",  x"95",  x"f1",  x"21",  x"03", -- 0740
         x"4b",  x"22",  x"c0",  x"f0",  x"21",  x"00",  x"00",  x"22", -- 0748
         x"c2",  x"f0",  x"3a",  x"6b",  x"f1",  x"d6",  x"0a",  x"32", -- 0750
         x"6f",  x"f1",  x"3a",  x"5b",  x"f1",  x"c6",  x"0a",  x"32", -- 0758
         x"5f",  x"f1",  x"21",  x"d5",  x"4a",  x"22",  x"b8",  x"f0", -- 0760
         x"21",  x"00",  x"00",  x"22",  x"ba",  x"f0",  x"0e",  x"64", -- 0768
         x"21",  x"b8",  x"f0",  x"3e",  x"04",  x"cd",  x"62",  x"48", -- 0770
         x"21",  x"c0",  x"f0",  x"3e",  x"0b",  x"cd",  x"62",  x"48", -- 0778
         x"cd",  x"9f",  x"1a",  x"79",  x"0f",  x"0f",  x"0f",  x"e6", -- 0780
         x"e0",  x"c2",  x"9a",  x"47",  x"3a",  x"6f",  x"f1",  x"3c", -- 0788
         x"32",  x"6f",  x"f1",  x"3a",  x"70",  x"f1",  x"3c",  x"32", -- 0790
         x"70",  x"f1",  x"0d",  x"c2",  x"70",  x"47",  x"21",  x"00", -- 0798
         x"00",  x"22",  x"7f",  x"f1",  x"cd",  x"2c",  x"24",  x"cd", -- 07A0
         x"9f",  x"1a",  x"c3",  x"85",  x"45",  x"3e",  x"ff",  x"32", -- 07A8
         x"b0",  x"f0",  x"32",  x"19",  x"f1",  x"21",  x"05",  x"4b", -- 07B0
         x"22",  x"c4",  x"f0",  x"21",  x"00",  x"00",  x"22",  x"c6", -- 07B8
         x"f0",  x"3a",  x"5f",  x"f1",  x"c6",  x"07",  x"32",  x"65", -- 07C0
         x"f1",  x"3a",  x"6f",  x"f1",  x"c6",  x"14",  x"32",  x"75", -- 07C8
         x"f1",  x"3e",  x"59",  x"32",  x"a6",  x"f1",  x"21",  x"bb", -- 07D0
         x"4a",  x"c3",  x"ac",  x"46",  x"21",  x"00",  x"00",  x"22", -- 07D8
         x"7b",  x"f1",  x"22",  x"7d",  x"f1",  x"21",  x"bc",  x"f0", -- 07E0
         x"3e",  x"00",  x"cd",  x"62",  x"48",  x"cd",  x"9f",  x"1a", -- 07E8
         x"d2",  x"e5",  x"47",  x"21",  x"00",  x"00",  x"22",  x"7b", -- 07F0
         x"f1",  x"22",  x"7d",  x"f1",  x"3e",  x"04",  x"32",  x"95", -- 07F8
         x"f1",  x"21",  x"e0",  x"f0",  x"22",  x"6b",  x"f1",  x"22", -- 0800
         x"6d",  x"f1",  x"3a",  x"6f",  x"f1",  x"fe",  x"8c",  x"da", -- 0808
         x"a1",  x"46",  x"3e",  x"ff",  x"32",  x"b3",  x"f0",  x"c3", -- 0810
         x"a1",  x"46",  x"af",  x"32",  x"19",  x"f1",  x"3e",  x"ff", -- 0818
         x"32",  x"b0",  x"f0",  x"c9",  x"c5",  x"d5",  x"e5",  x"f5", -- 0820
         x"21",  x"7b",  x"f1",  x"16",  x"00",  x"19",  x"eb",  x"21", -- 0828
         x"5b",  x"4b",  x"cd",  x"c6",  x"48",  x"d2",  x"53",  x"48", -- 0830
         x"21",  x"53",  x"4b",  x"cd",  x"c6",  x"48",  x"d2",  x"53", -- 0838
         x"48",  x"21",  x"15",  x"4b",  x"cd",  x"c6",  x"48",  x"d2", -- 0840
         x"53",  x"48",  x"21",  x"ec",  x"17",  x"cd",  x"c6",  x"48", -- 0848
         x"da",  x"79",  x"49",  x"23",  x"4e",  x"23",  x"7e",  x"12", -- 0850
         x"13",  x"0d",  x"c2",  x"55",  x"48",  x"f1",  x"e1",  x"d1", -- 0858
         x"c1",  x"c9",  x"32",  x"b2",  x"f0",  x"c5",  x"d5",  x"e5", -- 0860
         x"f5",  x"5e",  x"23",  x"56",  x"23",  x"06",  x"00",  x"4e", -- 0868
         x"eb",  x"09",  x"46",  x"eb",  x"79",  x"b7",  x"c2",  x"8f", -- 0870
         x"48",  x"78",  x"06",  x"00",  x"48",  x"cd",  x"f7",  x"48", -- 0878
         x"34",  x"34",  x"34",  x"34",  x"f1",  x"37",  x"3f",  x"e1", -- 0880
         x"d1",  x"c1",  x"c9",  x"35",  x"c3",  x"84",  x"48",  x"23", -- 0888
         x"7e",  x"b7",  x"c2",  x"8b",  x"48",  x"1b",  x"1b",  x"1b", -- 0890
         x"1a",  x"fe",  x"2e",  x"ca",  x"bb",  x"48",  x"fe",  x"2f", -- 0898
         x"ca",  x"b3",  x"48",  x"47",  x"13",  x"1a",  x"4f",  x"13", -- 08A0
         x"1a",  x"77",  x"13",  x"1a",  x"cd",  x"f7",  x"48",  x"2b", -- 08A8
         x"c3",  x"80",  x"48",  x"36",  x"00",  x"2b",  x"36",  x"00", -- 08B0
         x"c3",  x"84",  x"48",  x"36",  x"00",  x"2b",  x"36",  x"00", -- 08B8
         x"f1",  x"37",  x"e1",  x"d1",  x"c1",  x"c9",  x"c5",  x"d5", -- 08C0
         x"e5",  x"f5",  x"11",  x"06",  x"00",  x"be",  x"ca",  x"dd", -- 08C8
         x"48",  x"4f",  x"7e",  x"fe",  x"2f",  x"79",  x"ca",  x"e4", -- 08D0
         x"48",  x"19",  x"c3",  x"cd",  x"48",  x"f1",  x"37",  x"3f", -- 08D8
         x"d1",  x"d1",  x"c1",  x"c9",  x"f1",  x"37",  x"e1",  x"d1", -- 08E0
         x"c1",  x"c9",  x"85",  x"6f",  x"d0",  x"24",  x"c9",  x"af", -- 08E8
         x"02",  x"03",  x"1d",  x"c2",  x"f0",  x"48",  x"c9",  x"c5", -- 08F0
         x"d5",  x"e5",  x"f5",  x"21",  x"b2",  x"f0",  x"5e",  x"cd", -- 08F8
         x"24",  x"48",  x"1e",  x"0b",  x"21",  x"5b",  x"4b",  x"cd", -- 0900
         x"c6",  x"48",  x"d2",  x"2e",  x"49",  x"1e",  x"07",  x"21", -- 0908
         x"53",  x"4b",  x"cd",  x"c6",  x"48",  x"d2",  x"2e",  x"49", -- 0910
         x"1e",  x"09",  x"21",  x"15",  x"4b",  x"cd",  x"c6",  x"48", -- 0918
         x"d2",  x"2e",  x"49",  x"1e",  x"05",  x"21",  x"ec",  x"17", -- 0920
         x"cd",  x"c6",  x"48",  x"da",  x"79",  x"49",  x"23",  x"56", -- 0928
         x"23",  x"7e",  x"c5",  x"e5",  x"21",  x"7b",  x"f1",  x"f5", -- 0930
         x"3a",  x"b2",  x"f0",  x"cd",  x"ea",  x"48",  x"f1",  x"0e", -- 0938
         x"04",  x"be",  x"ca",  x"4f",  x"49",  x"23",  x"0d",  x"c2", -- 0940
         x"41",  x"49",  x"e1",  x"c1",  x"c3",  x"79",  x"49",  x"e1", -- 0948
         x"3a",  x"b2",  x"f0",  x"c6",  x"04",  x"91",  x"c1",  x"e5", -- 0950
         x"21",  x"5b",  x"f1",  x"cd",  x"ea",  x"48",  x"7e",  x"81", -- 0958
         x"77",  x"3e",  x"10",  x"cd",  x"ea",  x"48",  x"7e",  x"80", -- 0960
         x"77",  x"3e",  x"20",  x"cd",  x"ea",  x"48",  x"73",  x"e1", -- 0968
         x"15",  x"c2",  x"30",  x"49",  x"f1",  x"e1",  x"d1",  x"c1", -- 0970
         x"c9",  x"c3",  x"74",  x"49",  x"c5",  x"d5",  x"e5",  x"f5", -- 0978
         x"5e",  x"23",  x"56",  x"23",  x"4e",  x"23",  x"7e",  x"12", -- 0980
         x"23",  x"13",  x"0d",  x"c2",  x"86",  x"49",  x"f1",  x"e1", -- 0988
         x"d1",  x"c1",  x"c9",  x"91",  x"d0",  x"2f",  x"3c",  x"c9", -- 0990
         x"c5",  x"d5",  x"e5",  x"f5",  x"21",  x"be",  x"49",  x"0e", -- 0998
         x"06",  x"be",  x"ca",  x"b2",  x"49",  x"23",  x"23",  x"23", -- 09A0
         x"0d",  x"c2",  x"a1",  x"49",  x"f1",  x"37",  x"e1",  x"d1", -- 09A8
         x"c1",  x"c9",  x"23",  x"5e",  x"23",  x"56",  x"eb",  x"f1", -- 09B0
         x"37",  x"3f",  x"d1",  x"d1",  x"c1",  x"c9",  x"4a",  x"f2", -- 09B8
         x"46",  x"4c",  x"e4",  x"46",  x"59",  x"ad",  x"47",  x"42", -- 09C0
         x"ce",  x"46",  x"47",  x"b8",  x"46",  x"53",  x"a1",  x"46", -- 09C8
         x"b4",  x"f0",  x"18",  x"eb",  x"49",  x"00",  x"00",  x"6d", -- 09D0
         x"4a",  x"00",  x"00",  x"df",  x"4a",  x"00",  x"00",  x"f1", -- 09D8
         x"4a",  x"00",  x"00",  x"05",  x"4b",  x"00",  x"00",  x"0b", -- 09E0
         x"4b",  x"00",  x"00",  x"01",  x"00",  x"00",  x"04",  x"3c", -- 09E8
         x"04",  x"00",  x"04",  x"02",  x"fc",  x"00",  x"04",  x"31", -- 09F0
         x"00",  x"00",  x"04",  x"01",  x"00",  x"00",  x"03",  x"3c", -- 09F8
         x"04",  x"00",  x"03",  x"02",  x"fc",  x"00",  x"03",  x"31", -- 0A00
         x"00",  x"00",  x"03",  x"01",  x"00",  x"00",  x"02",  x"3c", -- 0A08
         x"04",  x"00",  x"02",  x"02",  x"fc",  x"00",  x"02",  x"31", -- 0A10
         x"00",  x"00",  x"02",  x"01",  x"00",  x"00",  x"01",  x"01", -- 0A18
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A20
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A28
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A30
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A38
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A40
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A48
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A50
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A58
         x"00",  x"00",  x"01",  x"1e",  x"00",  x"00",  x"01",  x"01", -- 0A60
         x"00",  x"00",  x"01",  x"1e",  x"2e",  x"46",  x"00",  x"00", -- 0A68
         x"08",  x"46",  x"2f",  x"34",  x"ff",  x"00",  x"07",  x"35", -- 0A70
         x"08",  x"00",  x"07",  x"36",  x"ff",  x"00",  x"07",  x"37", -- 0A78
         x"08",  x"00",  x"07",  x"34",  x"2f",  x"46",  x"fd",  x"00", -- 0A80
         x"09",  x"34",  x"fd",  x"00",  x"09",  x"46",  x"2f",  x"3b", -- 0A88
         x"00",  x"00",  x"04",  x"3b",  x"2f",  x"4a",  x"fe",  x"00", -- 0A90
         x"04",  x"46",  x"fa",  x"00",  x"04",  x"47",  x"04",  x"fb", -- 0A98
         x"04",  x"47",  x"0c",  x"fa",  x"04",  x"48",  x"06",  x"ff", -- 0AA0
         x"04",  x"48",  x"06",  x"01",  x"04",  x"48",  x"06",  x"05", -- 0AA8
         x"04",  x"49",  x"04",  x"06",  x"04",  x"49",  x"0e",  x"00", -- 0AB0
         x"06",  x"4a",  x"2e",  x"4a",  x"fe",  x"00",  x"04",  x"46", -- 0AB8
         x"f8",  x"00",  x"04",  x"38",  x"fb",  x"00",  x"08",  x"39", -- 0AC0
         x"10",  x"00",  x"0c",  x"3a",  x"f7",  x"00",  x"09",  x"38", -- 0AC8
         x"08",  x"00",  x"07",  x"46",  x"2e",  x"c3",  x"00",  x"00", -- 0AD0
         x"03",  x"c4",  x"00",  x"00",  x"03",  x"c3",  x"2f",  x"25", -- 0AD8
         x"00",  x"00",  x"06",  x"26",  x"00",  x"00",  x"06",  x"27", -- 0AE0
         x"00",  x"00",  x"06",  x"28",  x"00",  x"00",  x"06",  x"25", -- 0AE8
         x"2e",  x"1e",  x"fc",  x"00",  x"02",  x"1f",  x"fc",  x"00", -- 0AF0
         x"02",  x"20",  x"fc",  x"00",  x"02",  x"21",  x"fc",  x"00", -- 0AF8
         x"02",  x"1e",  x"2f",  x"1e",  x"2e",  x"4d",  x"00",  x"00", -- 0B00
         x"04",  x"4d",  x"2e",  x"03",  x"00",  x"00",  x"08",  x"04", -- 0B08
         x"00",  x"00",  x"08",  x"03",  x"2f",  x"31",  x"04",  x"b7", -- 0B10
         x"50",  x"7f",  x"7e",  x"1e",  x"04",  x"00",  x"40",  x"70", -- 0B18
         x"60",  x"1f",  x"04",  x"51",  x"41",  x"71",  x"61",  x"20", -- 0B20
         x"04",  x"00",  x"40",  x"52",  x"42",  x"21",  x"04",  x"51", -- 0B28
         x"41",  x"72",  x"62",  x"0d",  x"01",  x"4e",  x"00",  x"00", -- 0B30
         x"00",  x"0e",  x"01",  x"4f",  x"00",  x"00",  x"00",  x"0f", -- 0B38
         x"01",  x"5a",  x"00",  x"00",  x"00",  x"10",  x"01",  x"5b", -- 0B40
         x"00",  x"00",  x"00",  x"c0",  x"04",  x"00",  x"d8",  x"f8", -- 0B48
         x"e8",  x"2f",  x"2e",  x"c1",  x"04",  x"e8",  x"f8",  x"d8", -- 0B50
         x"00",  x"2f",  x"2e",  x"c2",  x"04",  x"f8",  x"e8",  x"00", -- 0B58
         x"d8",  x"2f",  x"2e",  x"5b",  x"f1",  x"40",  x"98",  x"98", -- 0B60
         x"a8",  x"a8",  x"98",  x"98",  x"a8",  x"a8",  x"90",  x"90", -- 0B68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"c0",  x"d0", -- 0B70
         x"c0",  x"d0",  x"10",  x"20",  x"10",  x"20",  x"40",  x"50", -- 0B78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0B88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"04",  x"04", -- 0B90
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B98
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"3e",  x"0d", -- 0BA0
         x"c3",  x"ad",  x"4b",  x"3e",  x"0b",  x"32",  x"0b",  x"f1", -- 0BA8
         x"3e",  x"01",  x"32",  x"ec",  x"f0",  x"cd",  x"af",  x"4d", -- 0BB0
         x"cd",  x"d5",  x"53",  x"cd",  x"9f",  x"1a",  x"af",  x"32", -- 0BB8
         x"19",  x"f1",  x"32",  x"b3",  x"f0",  x"32",  x"d1",  x"f0", -- 0BC0
         x"3e",  x"ff",  x"32",  x"b0",  x"f0",  x"3e",  x"53",  x"32", -- 0BC8
         x"a6",  x"f1",  x"cd",  x"9f",  x"1a",  x"cd",  x"16",  x"4e", -- 0BD0
         x"cd",  x"ec",  x"50",  x"3a",  x"a6",  x"f1",  x"fe",  x"59", -- 0BD8
         x"c2",  x"01",  x"4c",  x"3a",  x"ba",  x"f0",  x"fe",  x"14", -- 0BE0
         x"c2",  x"01",  x"4c",  x"21",  x"c4",  x"f0",  x"3e",  x"0a", -- 0BE8
         x"cd",  x"62",  x"48",  x"cd",  x"9f",  x"1a",  x"d2",  x"eb", -- 0BF0
         x"4b",  x"3e",  x"04",  x"32",  x"95",  x"f1",  x"c3",  x"4f", -- 0BF8
         x"4c",  x"3a",  x"b0",  x"f0",  x"b7",  x"ca",  x"1d",  x"4c", -- 0C00
         x"21",  x"b8",  x"f0",  x"3e",  x"04",  x"cd",  x"62",  x"48", -- 0C08
         x"d2",  x"1d",  x"4c",  x"af",  x"32",  x"b0",  x"f0",  x"32", -- 0C10
         x"19",  x"f1",  x"32",  x"a6",  x"f1",  x"3a",  x"6f",  x"f1", -- 0C18
         x"fe",  x"f0",  x"da",  x"3e",  x"4c",  x"3a",  x"d1",  x"f0", -- 0C20
         x"fe",  x"02",  x"d0",  x"3a",  x"6f",  x"f1",  x"c6",  x"04", -- 0C28
         x"32",  x"6f",  x"f1",  x"32",  x"71",  x"f1",  x"c6",  x"10", -- 0C30
         x"32",  x"70",  x"f1",  x"32",  x"72",  x"f1",  x"3a",  x"19", -- 0C38
         x"f1",  x"b7",  x"c2",  x"d2",  x"4b",  x"cd",  x"b6",  x"20", -- 0C40
         x"cd",  x"ea",  x"4c",  x"da",  x"d2",  x"4b",  x"e9",  x"cd", -- 0C48
         x"1a",  x"48",  x"3e",  x"53",  x"32",  x"a6",  x"f1",  x"21", -- 0C50
         x"6d",  x"4a",  x"22",  x"b8",  x"f0",  x"21",  x"00",  x"00", -- 0C58
         x"22",  x"ba",  x"f0",  x"c3",  x"d2",  x"4b",  x"3a",  x"a6", -- 0C60
         x"f1",  x"fe",  x"47",  x"ca",  x"d2",  x"4b",  x"cd",  x"1a", -- 0C68
         x"48",  x"3e",  x"47",  x"32",  x"a6",  x"f1",  x"21",  x"73", -- 0C70
         x"4a",  x"c3",  x"5a",  x"4c",  x"3a",  x"a6",  x"f1",  x"fe", -- 0C78
         x"42",  x"ca",  x"d2",  x"4b",  x"3a",  x"0b",  x"f1",  x"fe", -- 0C80
         x"0d",  x"ca",  x"d2",  x"4b",  x"cd",  x"1a",  x"48",  x"3e", -- 0C88
         x"42",  x"32",  x"a6",  x"f1",  x"21",  x"85",  x"4a",  x"c3", -- 0C90
         x"5a",  x"4c",  x"cd",  x"1a",  x"48",  x"3e",  x"4c",  x"32", -- 0C98
         x"a6",  x"f1",  x"21",  x"8f",  x"4a",  x"c3",  x"5a",  x"4c", -- 0CA0
         x"3e",  x"ff",  x"32",  x"b0",  x"f0",  x"32",  x"19",  x"f1", -- 0CA8
         x"3e",  x"4a",  x"32",  x"a6",  x"f1",  x"21",  x"95",  x"4a", -- 0CB0
         x"c3",  x"5a",  x"4c",  x"3e",  x"ff",  x"32",  x"b0",  x"f0", -- 0CB8
         x"32",  x"19",  x"f1",  x"21",  x"05",  x"4b",  x"22",  x"c4", -- 0CC0
         x"f0",  x"21",  x"00",  x"00",  x"22",  x"c6",  x"f0",  x"3a", -- 0CC8
         x"5f",  x"f1",  x"c6",  x"07",  x"32",  x"65",  x"f1",  x"3a", -- 0CD0
         x"6f",  x"f1",  x"c6",  x"14",  x"32",  x"75",  x"f1",  x"3e", -- 0CD8
         x"59",  x"32",  x"a6",  x"f1",  x"21",  x"bb",  x"4a",  x"c3", -- 0CE0
         x"5a",  x"4c",  x"c5",  x"d5",  x"e5",  x"f5",  x"21",  x"10", -- 0CE8
         x"4d",  x"0e",  x"06",  x"be",  x"ca",  x"04",  x"4d",  x"23", -- 0CF0
         x"23",  x"23",  x"0d",  x"c2",  x"f3",  x"4c",  x"f1",  x"37", -- 0CF8
         x"e1",  x"d1",  x"c1",  x"c9",  x"23",  x"5e",  x"23",  x"56", -- 0D00
         x"eb",  x"f1",  x"37",  x"3f",  x"d1",  x"d1",  x"c1",  x"c9", -- 0D08
         x"4a",  x"a8",  x"4c",  x"4c",  x"9a",  x"4c",  x"59",  x"bb", -- 0D10
         x"4c",  x"42",  x"7c",  x"4c",  x"47",  x"66",  x"4c",  x"53", -- 0D18
         x"4f",  x"4c",  x"b8",  x"f0",  x"04",  x"6d",  x"4a",  x"00", -- 0D20
         x"00",  x"5b",  x"f1",  x"40",  x"6b",  x"00",  x"c0",  x"c0", -- 0D28
         x"a8",  x"a8",  x"b8",  x"b8",  x"72",  x"72",  x"00",  x"00", -- 0D30
         x"00",  x"00",  x"00",  x"00",  x"f0",  x"00",  x"56",  x"66", -- 0D38
         x"10",  x"20",  x"10",  x"20",  x"d8",  x"e8",  x"00",  x"00", -- 0D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"43",  x"63", -- 0D48
         x"00",  x"00",  x"00",  x"00",  x"43",  x"63",  x"00",  x"00", -- 0D50
         x"00",  x"00",  x"00",  x"00",  x"05",  x"04",  x"05",  x"05", -- 0D58
         x"04",  x"04",  x"04",  x"04",  x"05",  x"05",  x"04",  x"04", -- 0D60
         x"04",  x"04",  x"04",  x"04",  x"5b",  x"f1",  x"40",  x"6c", -- 0D68
         x"00",  x"00",  x"00",  x"a8",  x"a8",  x"b8",  x"b8",  x"88", -- 0D70
         x"88",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"c0", -- 0D78
         x"00",  x"00",  x"00",  x"06",  x"16",  x"06",  x"16",  x"30", -- 0D80
         x"40",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0D88
         x"00",  x"43",  x"63",  x"00",  x"00",  x"00",  x"00",  x"43", -- 0D90
         x"63",  x"00",  x"00",  x"00",  x"00",  x"43",  x"63",  x"05", -- 0D98
         x"05",  x"05",  x"05",  x"05",  x"05",  x"05",  x"05",  x"05", -- 0DA0
         x"05",  x"05",  x"05",  x"05",  x"05",  x"05",  x"05",  x"3a", -- 0DA8
         x"0b",  x"f1",  x"fe",  x"0b",  x"c0",  x"21",  x"29",  x"4d", -- 0DB0
         x"cd",  x"7c",  x"49",  x"21",  x"22",  x"4d",  x"cd",  x"7c", -- 0DB8
         x"49",  x"cd",  x"d4",  x"4d",  x"cd",  x"ef",  x"4d",  x"21", -- 0DC0
         x"05",  x"4b",  x"22",  x"c4",  x"f0",  x"21",  x"00",  x"00", -- 0DC8
         x"22",  x"c6",  x"f0",  x"c9",  x"21",  x"22",  x"54",  x"22", -- 0DD0
         x"cc",  x"f0",  x"21",  x"00",  x"00",  x"22",  x"ce",  x"f0", -- 0DD8
         x"af",  x"32",  x"d0",  x"f0",  x"3e",  x"f0",  x"32",  x"6b", -- 0DE0
         x"f1",  x"3e",  x"6b",  x"32",  x"5b",  x"f1",  x"c9",  x"21", -- 0DE8
         x"22",  x"17",  x"22",  x"c8",  x"f0",  x"21",  x"00",  x"00", -- 0DF0
         x"22",  x"ca",  x"f0",  x"3e",  x"50",  x"32",  x"66",  x"f1", -- 0DF8
         x"3e",  x"d0",  x"32",  x"76",  x"f1",  x"3a",  x"0b",  x"f1", -- 0E00
         x"fe",  x"0b",  x"c8",  x"3e",  x"3c",  x"32",  x"66",  x"f1", -- 0E08
         x"3e",  x"ec",  x"32",  x"76",  x"f1",  x"c9",  x"3a",  x"0b", -- 0E10
         x"f1",  x"fe",  x"0b",  x"c0",  x"21",  x"cc",  x"f0",  x"af", -- 0E18
         x"cd",  x"62",  x"48",  x"3a",  x"d0",  x"f0",  x"e6",  x"c0", -- 0E20
         x"ca",  x"37",  x"4e",  x"3a",  x"d0",  x"f0",  x"3d",  x"32", -- 0E28
         x"d0",  x"f0",  x"e6",  x"c0",  x"cc",  x"d4",  x"4d",  x"3a", -- 0E30
         x"d0",  x"f0",  x"b7",  x"c2",  x"57",  x"4e",  x"3a",  x"6b", -- 0E38
         x"f1",  x"fe",  x"68",  x"d2",  x"82",  x"4e",  x"21",  x"2c", -- 0E40
         x"54",  x"22",  x"cc",  x"f0",  x"21",  x"00",  x"00",  x"22", -- 0E48
         x"ce",  x"f0",  x"3e",  x"01",  x"32",  x"d0",  x"f0",  x"fe", -- 0E50
         x"01",  x"c2",  x"75",  x"4e",  x"3a",  x"5b",  x"f1",  x"fe", -- 0E58
         x"b8",  x"da",  x"82",  x"4e",  x"21",  x"22",  x"54",  x"22", -- 0E60
         x"cc",  x"f0",  x"21",  x"00",  x"00",  x"22",  x"ce",  x"f0", -- 0E68
         x"3e",  x"02",  x"32",  x"d0",  x"f0",  x"3a",  x"6b",  x"f1", -- 0E70
         x"fe",  x"08",  x"d2",  x"82",  x"4e",  x"3e",  x"ee",  x"32", -- 0E78
         x"d0",  x"f0",  x"3a",  x"d0",  x"f0",  x"fe",  x"01",  x"c2", -- 0E80
         x"a4",  x"4e",  x"3a",  x"5d",  x"f1",  x"4f",  x"3a",  x"5b", -- 0E88
         x"f1",  x"cd",  x"93",  x"49",  x"fe",  x"04",  x"d2",  x"a4", -- 0E90
         x"4e",  x"3a",  x"5d",  x"f1",  x"c6",  x"0a",  x"32",  x"5d", -- 0E98
         x"f1",  x"32",  x"5e",  x"f1",  x"3a",  x"b3",  x"f0",  x"fe", -- 0EA0
         x"04",  x"ca",  x"79",  x"50",  x"fe",  x"05",  x"d2",  x"7f", -- 0EA8
         x"50",  x"3a",  x"5f",  x"f1",  x"fe",  x"80",  x"da",  x"e9", -- 0EB0
         x"4e",  x"3a",  x"6f",  x"f1",  x"c6",  x"20",  x"d6",  x"8c", -- 0EB8
         x"da",  x"e9",  x"4e",  x"fe",  x"0a",  x"d2",  x"da",  x"4e", -- 0EC0
         x"3a",  x"6f",  x"f1",  x"d6",  x"0c",  x"6f",  x"c6",  x"10", -- 0EC8
         x"67",  x"22",  x"6f",  x"f1",  x"22",  x"71",  x"f1",  x"c3", -- 0ED0
         x"e9",  x"4e",  x"d6",  x"20",  x"fe",  x"08",  x"d2",  x"e9", -- 0ED8
         x"4e",  x"3a",  x"6f",  x"f1",  x"c6",  x"06",  x"c3",  x"cd", -- 0EE0
         x"4e",  x"3a",  x"6f",  x"f1",  x"d6",  x"04",  x"4f",  x"3a", -- 0EE8
         x"6d",  x"f1",  x"cd",  x"93",  x"49",  x"fe",  x"0a",  x"d2", -- 0EF0
         x"32",  x"4f",  x"3a",  x"a6",  x"f1",  x"fe",  x"53",  x"ca", -- 0EF8
         x"09",  x"4f",  x"3a",  x"ba",  x"f0",  x"b7",  x"c2",  x"32", -- 0F00
         x"4f",  x"3a",  x"5d",  x"f1",  x"d6",  x"01",  x"fe",  x"70", -- 0F08
         x"da",  x"24",  x"4f",  x"32",  x"5d",  x"f1",  x"32",  x"5e", -- 0F10
         x"f1",  x"3e",  x"01",  x"32",  x"b3",  x"f0",  x"cd",  x"d5", -- 0F18
         x"50",  x"c3",  x"32",  x"4f",  x"3a",  x"b3",  x"f0",  x"3d", -- 0F20
         x"c2",  x"32",  x"4f",  x"af",  x"32",  x"19",  x"f1",  x"32", -- 0F28
         x"b3",  x"f0",  x"3a",  x"6f",  x"f1",  x"d6",  x"04",  x"4f", -- 0F30
         x"3a",  x"73",  x"f1",  x"cd",  x"93",  x"49",  x"fe",  x"0a", -- 0F38
         x"d2",  x"81",  x"4f",  x"3a",  x"a6",  x"f1",  x"fe",  x"53", -- 0F40
         x"ca",  x"52",  x"4f",  x"3a",  x"ba",  x"f0",  x"b7",  x"c2", -- 0F48
         x"81",  x"4f",  x"3a",  x"63",  x"f1",  x"c6",  x"01",  x"fe", -- 0F50
         x"c0",  x"d2",  x"6d",  x"4f",  x"32",  x"63",  x"f1",  x"32", -- 0F58
         x"64",  x"f1",  x"3e",  x"02",  x"32",  x"b3",  x"f0",  x"cd", -- 0F60
         x"d5",  x"50",  x"c3",  x"81",  x"4f",  x"3e",  x"02",  x"32", -- 0F68
         x"d1",  x"f0",  x"3a",  x"b3",  x"f0",  x"fe",  x"02",  x"c2", -- 0F70
         x"81",  x"4f",  x"af",  x"32",  x"19",  x"f1",  x"32",  x"b3", -- 0F78
         x"f0",  x"3a",  x"6f",  x"f1",  x"4f",  x"3a",  x"6b",  x"f1", -- 0F80
         x"cd",  x"93",  x"49",  x"fe",  x"0a",  x"d2",  x"cf",  x"4f", -- 0F88
         x"3a",  x"d0",  x"f0",  x"3d",  x"ca",  x"cf",  x"4f",  x"3a", -- 0F90
         x"5f",  x"f1",  x"c6",  x"12",  x"4f",  x"3a",  x"5b",  x"f1", -- 0F98
         x"cd",  x"93",  x"49",  x"fe",  x"05",  x"d2",  x"cf",  x"4f", -- 0FA0
         x"21",  x"36",  x"54",  x"22",  x"cc",  x"f0",  x"3e",  x"ff", -- 0FA8
         x"32",  x"19",  x"f1",  x"32",  x"b0",  x"f0",  x"3e",  x"03", -- 0FB0
         x"32",  x"b3",  x"f0",  x"3e",  x"4c",  x"32",  x"a6",  x"f1", -- 0FB8
         x"21",  x"9c",  x"54",  x"22",  x"b8",  x"f0",  x"21",  x"00", -- 0FC0
         x"00",  x"22",  x"ba",  x"f0",  x"c3",  x"17",  x"50",  x"3a", -- 0FC8
         x"b3",  x"f0",  x"fe",  x"03",  x"c2",  x"ec",  x"4f",  x"3a", -- 0FD0
         x"ba",  x"f0",  x"b7",  x"c2",  x"ec",  x"4f",  x"cd",  x"2c", -- 0FD8
         x"24",  x"af",  x"32",  x"19",  x"f1",  x"32",  x"b3",  x"f0", -- 0FE0
         x"2f",  x"32",  x"b0",  x"f0",  x"3a",  x"b3",  x"f0",  x"3d", -- 0FE8
         x"c2",  x"09",  x"50",  x"3a",  x"5d",  x"f1",  x"d6",  x"1a", -- 0FF0
         x"32",  x"5f",  x"f1",  x"32",  x"60",  x"f1",  x"c6",  x"10", -- 0FF8
         x"32",  x"61",  x"f1",  x"32",  x"62",  x"f1",  x"c3",  x"17", -- 1000
         x"50",  x"3a",  x"b3",  x"f0",  x"fe",  x"02",  x"c2",  x"17", -- 1008
         x"50",  x"3a",  x"63",  x"f1",  x"c3",  x"f6",  x"4f",  x"3a", -- 1010
         x"76",  x"f1",  x"4f",  x"3a",  x"6f",  x"f1",  x"cd",  x"93", -- 1018
         x"49",  x"fe",  x"08",  x"d2",  x"5a",  x"50",  x"3a",  x"66", -- 1020
         x"f1",  x"4f",  x"3a",  x"5f",  x"f1",  x"cd",  x"93",  x"49", -- 1028
         x"fe",  x"08",  x"d2",  x"5a",  x"50",  x"3a",  x"a6",  x"f1", -- 1030
         x"fe",  x"4c",  x"ca",  x"5a",  x"50",  x"fe",  x"59",  x"c2", -- 1038
         x"4d",  x"50",  x"3a",  x"66",  x"f1",  x"d6",  x"10",  x"32", -- 1040
         x"66",  x"f1",  x"c3",  x"5a",  x"50",  x"3e",  x"50",  x"32", -- 1048
         x"66",  x"f1",  x"3e",  x"04",  x"32",  x"b3",  x"f0",  x"cd", -- 1050
         x"d5",  x"50",  x"21",  x"c8",  x"f0",  x"3e",  x"0b",  x"cd", -- 1058
         x"62",  x"48",  x"3a",  x"76",  x"f1",  x"fe",  x"24",  x"d2", -- 1060
         x"78",  x"50",  x"cd",  x"ef",  x"4d",  x"3a",  x"b3",  x"f0", -- 1068
         x"fe",  x"04",  x"c0",  x"3e",  x"05",  x"32",  x"b3",  x"f0", -- 1070
         x"c9",  x"cd",  x"b2",  x"50",  x"c3",  x"5a",  x"50",  x"3a", -- 1078
         x"b3",  x"f0",  x"fe",  x"06",  x"ca",  x"a0",  x"50",  x"21", -- 1080
         x"a2",  x"54",  x"22",  x"b8",  x"f0",  x"21",  x"00",  x"00", -- 1088
         x"22",  x"ba",  x"f0",  x"3e",  x"06",  x"32",  x"b3",  x"f0", -- 1090
         x"3e",  x"50",  x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f", -- 1098
         x"3a",  x"6f",  x"f1",  x"fe",  x"10",  x"da",  x"ab",  x"50", -- 10A0
         x"c3",  x"5a",  x"50",  x"f1",  x"cd",  x"2c",  x"24",  x"c3", -- 10A8
         x"b5",  x"4b",  x"3a",  x"76",  x"f1",  x"c6",  x"09",  x"6f", -- 10B0
         x"c6",  x"10",  x"67",  x"22",  x"6f",  x"f1",  x"22",  x"71", -- 10B8
         x"f1",  x"3a",  x"66",  x"f1",  x"c6",  x"04",  x"32",  x"5f", -- 10C0
         x"f1",  x"32",  x"60",  x"f1",  x"c6",  x"10",  x"32",  x"61", -- 10C8
         x"f1",  x"32",  x"62",  x"f1",  x"c9",  x"3e",  x"ff",  x"32", -- 10D0
         x"19",  x"f1",  x"3e",  x"53",  x"32",  x"a6",  x"f1",  x"21", -- 10D8
         x"6d",  x"4a",  x"22",  x"b8",  x"f0",  x"21",  x"00",  x"00", -- 10E0
         x"22",  x"ba",  x"f0",  x"c9",  x"3a",  x"0b",  x"f1",  x"fe", -- 10E8
         x"0d",  x"c0",  x"21",  x"bc",  x"f0",  x"af",  x"cd",  x"62", -- 10F0
         x"48",  x"da",  x"14",  x"52",  x"3a",  x"8f",  x"f1",  x"fe", -- 10F8
         x"04",  x"ca",  x"e3",  x"51",  x"3a",  x"72",  x"f1",  x"57", -- 1100
         x"3a",  x"6b",  x"f1",  x"47",  x"3a",  x"62",  x"f1",  x"5f", -- 1108
         x"3a",  x"5b",  x"f1",  x"4f",  x"7b",  x"cd",  x"93",  x"49", -- 1110
         x"5f",  x"48",  x"7a",  x"cd",  x"93",  x"49",  x"83",  x"da", -- 1118
         x"e3",  x"51",  x"fe",  x"10",  x"d2",  x"7c",  x"51",  x"4f", -- 1120
         x"3a",  x"a6",  x"f1",  x"fe",  x"59",  x"79",  x"ca",  x"5a", -- 1128
         x"51",  x"fe",  x"08",  x"d2",  x"7c",  x"51",  x"21",  x"04", -- 1130
         x"04",  x"22",  x"8f",  x"f1",  x"22",  x"91",  x"f1",  x"af", -- 1138
         x"32",  x"b0",  x"f0",  x"21",  x"df",  x"4a",  x"22",  x"bc", -- 1140
         x"f0",  x"21",  x"00",  x"00",  x"22",  x"be",  x"f0",  x"3e", -- 1148
         x"45",  x"32",  x"a6",  x"f1",  x"cd",  x"e3",  x"0f",  x"c3", -- 1150
         x"e3",  x"51",  x"3a",  x"bb",  x"f0",  x"2f",  x"e6",  x"03", -- 1158
         x"87",  x"4f",  x"06",  x"00",  x"21",  x"74",  x"51",  x"09", -- 1160
         x"7e",  x"32",  x"6b",  x"f1",  x"23",  x"7e",  x"32",  x"5b", -- 1168
         x"f1",  x"c3",  x"e3",  x"51",  x"c0",  x"6c",  x"90",  x"a2", -- 1170
         x"a8",  x"a2",  x"a8",  x"a2",  x"3a",  x"bb",  x"f0",  x"fe", -- 1178
         x"08",  x"c2",  x"e3",  x"51",  x"3a",  x"6f",  x"f1",  x"4f", -- 1180
         x"3a",  x"5f",  x"f1",  x"47",  x"3a",  x"6b",  x"f1",  x"5f", -- 1188
         x"3a",  x"5b",  x"f1",  x"81",  x"80",  x"83",  x"fe",  x"d2", -- 1190
         x"d2",  x"e3",  x"51",  x"3a",  x"8f",  x"f1",  x"fe",  x"04", -- 1198
         x"ca",  x"e3",  x"51",  x"3a",  x"6b",  x"f1",  x"5f",  x"3a", -- 11A0
         x"72",  x"f1",  x"57",  x"bb",  x"da",  x"b4",  x"51",  x"7b", -- 11A8
         x"c6",  x"04",  x"5f",  x"7a",  x"83",  x"1f",  x"83",  x"1f", -- 11B0
         x"83",  x"1f",  x"47",  x"32",  x"6b",  x"f1",  x"3a",  x"5b", -- 11B8
         x"f1",  x"4f",  x"3a",  x"62",  x"f1",  x"5f",  x"b9",  x"d2", -- 11C0
         x"cf",  x"51",  x"79",  x"d6",  x"02",  x"4f",  x"7b",  x"81", -- 11C8
         x"1f",  x"81",  x"1f",  x"81",  x"1f",  x"4f",  x"fe",  x"18", -- 11D0
         x"da",  x"e3",  x"51",  x"fe",  x"e0",  x"d2",  x"e3",  x"51", -- 11D8
         x"32",  x"5b",  x"f1",  x"3a",  x"76",  x"f1",  x"fe",  x"06", -- 11E0
         x"d2",  x"1b",  x"52",  x"cd",  x"ef",  x"4d",  x"af",  x"32", -- 11E8
         x"d2",  x"f0",  x"3a",  x"b3",  x"f0",  x"fe",  x"02",  x"c2", -- 11F0
         x"1b",  x"52",  x"21",  x"04",  x"04",  x"22",  x"8f",  x"f1", -- 11F8
         x"22",  x"91",  x"f1",  x"3e",  x"50",  x"32",  x"a6",  x"f1", -- 1200
         x"cd",  x"e3",  x"0f",  x"3e",  x"64",  x"cd",  x"9f",  x"1a", -- 1208
         x"3d",  x"c2",  x"0d",  x"52",  x"cd",  x"2c",  x"24",  x"f1", -- 1210
         x"c3",  x"b5",  x"4b",  x"21",  x"c8",  x"f0",  x"3e",  x"0b", -- 1218
         x"cd",  x"62",  x"48",  x"16",  x"00",  x"3a",  x"6f",  x"f1", -- 1220
         x"4f",  x"3a",  x"5f",  x"f1",  x"47",  x"21",  x"68",  x"54", -- 1228
         x"3a",  x"d2",  x"f0",  x"b7",  x"ca",  x"3f",  x"52",  x"16", -- 1230
         x"ff",  x"01",  x"10",  x"10",  x"21",  x"82",  x"54",  x"3a", -- 1238
         x"76",  x"f1",  x"22",  x"c8",  x"f0",  x"21",  x"22",  x"17", -- 1240
         x"3a",  x"66",  x"f1",  x"4f",  x"7a",  x"b7",  x"79",  x"ca", -- 1248
         x"5c",  x"52",  x"b8",  x"d2",  x"60",  x"52",  x"22",  x"c8", -- 1250
         x"f0",  x"c3",  x"60",  x"52",  x"b8",  x"d2",  x"56",  x"52", -- 1258
         x"3a",  x"b3",  x"f0",  x"fe",  x"02",  x"ca",  x"8b",  x"53", -- 1260
         x"b7",  x"ca",  x"c3",  x"52",  x"3a",  x"6d",  x"f1",  x"6f", -- 1268
         x"c6",  x"10",  x"67",  x"22",  x"6f",  x"f1",  x"22",  x"71", -- 1270
         x"f1",  x"3a",  x"5d",  x"f1",  x"d6",  x"1a",  x"6f",  x"67", -- 1278
         x"22",  x"5f",  x"f1",  x"c6",  x"10",  x"67",  x"6f",  x"22", -- 1280
         x"61",  x"f1",  x"21",  x"d3",  x"f0",  x"3a",  x"5d",  x"f1", -- 1288
         x"86",  x"23",  x"4f",  x"7e",  x"b7",  x"79",  x"23",  x"ca", -- 1290
         x"a1",  x"52",  x"be",  x"da",  x"be",  x"52",  x"c3",  x"a5", -- 1298
         x"52",  x"be",  x"d2",  x"be",  x"52",  x"3e",  x"00",  x"32", -- 12A0
         x"b3",  x"f0",  x"3a",  x"d1",  x"f0",  x"3c",  x"fe",  x"03", -- 12A8
         x"c2",  x"b5",  x"52",  x"3e",  x"04",  x"32",  x"d1",  x"f0", -- 12B0
         x"cd",  x"8f",  x"53",  x"c3",  x"c3",  x"52",  x"69",  x"61", -- 12B8
         x"22",  x"5d",  x"f1",  x"3a",  x"6f",  x"f1",  x"0e",  x"38", -- 12C0
         x"cd",  x"93",  x"49",  x"5f",  x"3a",  x"5f",  x"f1",  x"0e", -- 12C8
         x"70",  x"cd",  x"93",  x"49",  x"83",  x"da",  x"33",  x"53", -- 12D0
         x"fe",  x"10",  x"d2",  x"33",  x"53",  x"21",  x"04",  x"04", -- 12D8
         x"22",  x"8f",  x"f1",  x"22",  x"91",  x"f1",  x"3e",  x"32", -- 12E0
         x"cd",  x"9f",  x"1a",  x"f5",  x"21",  x"c8",  x"f0",  x"3e", -- 12E8
         x"0b",  x"cd",  x"62",  x"48",  x"21",  x"bc",  x"f0",  x"af", -- 12F0
         x"cd",  x"62",  x"48",  x"f1",  x"3d",  x"c2",  x"e8",  x"52", -- 12F8
         x"21",  x"05",  x"05",  x"22",  x"8f",  x"f1",  x"22",  x"91", -- 1300
         x"f1",  x"3a",  x"ca",  x"f0",  x"0f",  x"0f",  x"0f",  x"01", -- 1308
         x"38",  x"46",  x"da",  x"18",  x"53",  x"01",  x"a8",  x"56", -- 1310
         x"68",  x"78",  x"c6",  x"10",  x"67",  x"22",  x"6f",  x"f1", -- 1318
         x"22",  x"71",  x"f1",  x"69",  x"61",  x"22",  x"5f",  x"f1", -- 1320
         x"79",  x"c6",  x"10",  x"6f",  x"67",  x"22",  x"61",  x"f1", -- 1328
         x"cd",  x"8f",  x"53",  x"3a",  x"6f",  x"f1",  x"d6",  x"04", -- 1330
         x"4f",  x"3a",  x"6d",  x"f1",  x"cd",  x"93",  x"49",  x"fe", -- 1338
         x"0a",  x"d2",  x"49",  x"53",  x"3e",  x"01",  x"32",  x"b3", -- 1340
         x"f0",  x"3a",  x"76",  x"f1",  x"4f",  x"3a",  x"6f",  x"f1", -- 1348
         x"cd",  x"93",  x"49",  x"5f",  x"3a",  x"66",  x"f1",  x"4f", -- 1350
         x"3a",  x"5f",  x"f1",  x"cd",  x"93",  x"49",  x"83",  x"da", -- 1358
         x"8a",  x"53",  x"fe",  x"0b",  x"d2",  x"8a",  x"53",  x"3e", -- 1360
         x"01",  x"32",  x"d2",  x"f0",  x"3a",  x"a6",  x"f1",  x"fe", -- 1368
         x"4c",  x"ca",  x"8a",  x"53",  x"fe",  x"59",  x"ca",  x"82", -- 1370
         x"53",  x"3e",  x"02",  x"32",  x"b3",  x"f0",  x"cd",  x"d5", -- 1378
         x"50",  x"c9",  x"3a",  x"66",  x"f1",  x"d6",  x"10",  x"32", -- 1380
         x"66",  x"f1",  x"c9",  x"cd",  x"b2",  x"50",  x"c9",  x"2a", -- 1388
         x"5d",  x"f1",  x"22",  x"69",  x"f1",  x"2a",  x"6d",  x"f1", -- 1390
         x"22",  x"79",  x"f1",  x"3a",  x"5f",  x"f1",  x"fe",  x"60", -- 1398
         x"d2",  x"a8",  x"53",  x"3e",  x"03",  x"32",  x"d1",  x"f0", -- 13A0
         x"3a",  x"d1",  x"f0",  x"4f",  x"87",  x"87",  x"81",  x"4f", -- 13A8
         x"06",  x"00",  x"21",  x"09",  x"54",  x"09",  x"7e",  x"32", -- 13B0
         x"6d",  x"f1",  x"c6",  x"10",  x"32",  x"6e",  x"f1",  x"23", -- 13B8
         x"7e",  x"32",  x"5d",  x"f1",  x"32",  x"5e",  x"f1",  x"23", -- 13C0
         x"7e",  x"32",  x"d3",  x"f0",  x"23",  x"5e",  x"23",  x"56", -- 13C8
         x"eb",  x"22",  x"d4",  x"f0",  x"c9",  x"3a",  x"0b",  x"f1", -- 13D0
         x"fe",  x"0d",  x"c0",  x"21",  x"6c",  x"4d",  x"cd",  x"7c", -- 13D8
         x"49",  x"af",  x"32",  x"d2",  x"f0",  x"32",  x"d1",  x"f0", -- 13E0
         x"67",  x"6f",  x"22",  x"c6",  x"f0",  x"22",  x"ba",  x"f0", -- 13E8
         x"22",  x"be",  x"f0",  x"21",  x"6d",  x"4a",  x"22",  x"b8", -- 13F0
         x"f0",  x"21",  x"05",  x"4b",  x"22",  x"c4",  x"f0",  x"21", -- 13F8
         x"b4",  x"54",  x"22",  x"bc",  x"f0",  x"cd",  x"8f",  x"53", -- 1400
         x"c9",  x"18",  x"c0",  x"ff",  x"00",  x"88",  x"68",  x"c0", -- 1408
         x"ff",  x"00",  x"88",  x"e0",  x"88",  x"01",  x"ff",  x"c0", -- 1410
         x"e0",  x"50",  x"01",  x"ff",  x"c0",  x"68",  x"c0",  x"ff", -- 1418
         x"00",  x"88",  x"06",  x"fc",  x"00",  x"01",  x"07",  x"fc", -- 1420
         x"00",  x"01",  x"06",  x"2f",  x"06",  x"ff",  x"04",  x"01", -- 1428
         x"07",  x"ff",  x"04",  x"01",  x"06",  x"2f",  x"06",  x"fd", -- 1430
         x"fe",  x"01",  x"07",  x"fd",  x"fe",  x"01",  x"06",  x"fd", -- 1438
         x"fe",  x"01",  x"07",  x"fd",  x"fe",  x"01",  x"06",  x"fd", -- 1440
         x"fe",  x"01",  x"07",  x"fd",  x"fe",  x"01",  x"06",  x"fd", -- 1448
         x"02",  x"01",  x"07",  x"fd",  x"02",  x"01",  x"06",  x"fd", -- 1450
         x"02",  x"01",  x"07",  x"fd",  x"02",  x"01",  x"06",  x"fd", -- 1458
         x"02",  x"01",  x"07",  x"fd",  x"02",  x"01",  x"06",  x"2f", -- 1460
         x"0d",  x"fd",  x"05",  x"02",  x"0e",  x"fd",  x"05",  x"02", -- 1468
         x"0f",  x"fd",  x"04",  x"02",  x"10",  x"fd",  x"05",  x"02", -- 1470
         x"0f",  x"fd",  x"05",  x"02",  x"0e",  x"fd",  x"06",  x"02", -- 1478
         x"0d",  x"2f",  x"0d",  x"fd",  x"fb",  x"02",  x"0e",  x"fd", -- 1480
         x"fb",  x"02",  x"0f",  x"fd",  x"fb",  x"02",  x"10",  x"fd", -- 1488
         x"fb",  x"02",  x"0f",  x"fd",  x"fb",  x"02",  x"0e",  x"fd", -- 1490
         x"fb",  x"02",  x"0d",  x"2f",  x"3b",  x"00",  x"00",  x"40", -- 1498
         x"3b",  x"2f",  x"46",  x"fd",  x"08",  x"05",  x"c0",  x"fd", -- 14A0
         x"08",  x"05",  x"c1",  x"fd",  x"08",  x"05",  x"c2",  x"fd", -- 14A8
         x"08",  x"05",  x"46",  x"2f",  x"25",  x"02",  x"00",  x"04", -- 14B0
         x"26",  x"00",  x"fe",  x"04",  x"25",  x"fe",  x"00",  x"04", -- 14B8
         x"26",  x"00",  x"02",  x"04",  x"25",  x"2f",  x"d3",  x"00", -- 14C0
         x"c9",  x"c1",  x"c3",  x"00",  x"00",  x"32",  x"00",  x"00", -- 14C8
         x"c9",  x"21",  x"00",  x"00",  x"c9",  x"21",  x"00",  x"00", -- 14D0
         x"c9",  x"32",  x"88",  x"f1",  x"32",  x"78",  x"f1",  x"c9", -- 14D8
         x"c6",  x"03",  x"c9",  x"c6",  x"fd",  x"c9",  x"fe",  x"bf", -- 14E0
         x"c9",  x"fe",  x"a7",  x"c9",  x"fe",  x"bf",  x"c9",  x"46", -- 14E8
         x"00",  x"00",  x"00",  x"46",  x"2f",  x"db",  x"d2",  x"e6", -- 14F0
         x"80",  x"ca",  x"2f",  x"f0",  x"3a",  x"f2",  x"f0",  x"b7", -- 14F8
         x"ca",  x"44",  x"f0",  x"3a",  x"ec",  x"f0",  x"b7",  x"c2", -- 1500
         x"59",  x"f0",  x"11",  x"1b",  x"f1",  x"21",  x"4e",  x"f0", -- 1508
         x"06",  x"40",  x"1a",  x"d3",  x"40",  x"13",  x"34",  x"05", -- 1510
         x"c2",  x"4c",  x"f0",  x"cd",  x"1b",  x"10",  x"c9",  x"cd", -- 1518
         x"a9",  x"14",  x"06",  x"1a",  x"11",  x"89",  x"f0",  x"21", -- 1520
         x"48",  x"15",  x"22",  x"68",  x"f0",  x"2a",  x"48",  x"15", -- 1528
         x"1a",  x"77",  x"05",  x"2a",  x"68",  x"f0",  x"23",  x"23", -- 1530
         x"13",  x"c2",  x"64",  x"f0",  x"3e",  x"00",  x"d3",  x"bd", -- 1538
         x"3e",  x"00",  x"d3",  x"bc",  x"cd",  x"b2",  x"14",  x"af", -- 1540
         x"32",  x"ec",  x"f0",  x"cd",  x"1b",  x"10",  x"c9",  x"ff", -- 1548
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1550
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1558
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1560
         x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1568
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 1570
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1578
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1580
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1588
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1590
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1598
         x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00",  x"00", -- 15A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 15A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 15B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 15B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 15C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 15C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"fe", -- 15D0
         x"02",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 15D8
         x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 15F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1600
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1608
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1610
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1618
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1620
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1628
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1630
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1638
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1640
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1648
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1650
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1658
         x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1660
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 1668
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1670
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1678
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1680
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1688
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1690
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1698
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 16F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1700
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1708
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1710
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1718
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1720
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1728
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1730
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1738
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1740
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1748
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1750
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1758
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1760
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1768
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1770
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1778
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1780
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1788
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1790
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1798
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 17F8
         x"00",  x"a9",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1810
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1828
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1838
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1848
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1850
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1868
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1878
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1880
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1888
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1890
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1898
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18F8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1900
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1908
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1910
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1918
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1920
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1928
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1930
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1938
         x"15",  x"15",  x"15",  x"5d",  x"2f",  x"22",  x"20",  x"17", -- 1940
         x"15",  x"15",  x"15",  x"13",  x"21",  x"22",  x"22",  x"20", -- 1948
         x"15",  x"13",  x"15",  x"21",  x"39",  x"15",  x"15",  x"15", -- 1950
         x"5d",  x"15",  x"15",  x"21",  x"22",  x"22",  x"20",  x"15", -- 1958
         x"15",  x"15",  x"15",  x"14",  x"54",  x"53",  x"2c",  x"4d", -- 1960
         x"16",  x"5c",  x"14",  x"13",  x"58",  x"52",  x"51",  x"2c", -- 1968
         x"14",  x"15",  x"15",  x"14",  x"54",  x"39",  x"17",  x"15", -- 1970
         x"15",  x"13",  x"15",  x"58",  x"54",  x"53",  x"15",  x"15", -- 1978
         x"12",  x"5c",  x"14",  x"58",  x"52",  x"51",  x"11",  x"0b", -- 1980
         x"10",  x"4d",  x"14",  x"15",  x"58",  x"54",  x"53",  x"11", -- 1988
         x"12",  x"5c",  x"14",  x"58",  x"52",  x"51",  x"14",  x"17", -- 1990
         x"11",  x"12",  x"14",  x"15",  x"52",  x"51",  x"2c",  x"4d", -- 1998
         x"0b",  x"12",  x"4d",  x"11",  x"54",  x"53",  x"0b",  x"0b", -- 19A0
         x"0b",  x"0b",  x"12",  x"4d",  x"11",  x"52",  x"51",  x"0b", -- 19A8
         x"10",  x"11",  x"12",  x"4d",  x"54",  x"53",  x"4d",  x"11", -- 19B0
         x"0b",  x"0b",  x"10",  x"4d",  x"54",  x"53",  x"11",  x"0b", -- 19B8
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b", -- 19C0
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23", -- 19C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"52",  x"51",  x"23",  x"0b", -- 19D0
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b", -- 19D8
         x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b", -- 19E0
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23", -- 19E8
         x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"0b",  x"0b", -- 19F0
         x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"23",  x"0b", -- 19F8
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b", -- 1A00
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"38",  x"29", -- 1A08
         x"30",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b", -- 1A10
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b", -- 1A18
         x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"0b",  x"0b", -- 1A20
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"52",  x"39",  x"4d", -- 1A28
         x"28",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"29",  x"30", -- 1A30
         x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"0b",  x"0b", -- 1A38
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"1b",  x"c1", -- 1A40
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23", -- 1A48
         x"c0",  x"c1",  x"0b",  x"0b",  x"52",  x"51",  x"4d",  x"28", -- 1A50
         x"0b",  x"0b",  x"0b",  x"0b",  x"52",  x"51",  x"23",  x"0b", -- 1A58
         x"2a",  x"c1",  x"0b",  x"2a",  x"54",  x"53",  x"04",  x"04", -- 1A60
         x"c1",  x"0b",  x"2a",  x"1f",  x"c0",  x"52",  x"51",  x"c1", -- 1A68
         x"04",  x"04",  x"1f",  x"2a",  x"54",  x"53",  x"c0",  x"c1", -- 1A70
         x"0b",  x"2a",  x"c1",  x"c0",  x"54",  x"53",  x"1f",  x"0b", -- 1A78
         x"04",  x"04",  x"1b",  x"26",  x"52",  x"51",  x"27",  x"04", -- 1A80
         x"04",  x"1b",  x"04",  x"1c",  x"26",  x"54",  x"53",  x"27", -- 1A88
         x"04",  x"04",  x"1c",  x"26",  x"52",  x"51",  x"27",  x"04", -- 1A90
         x"1b",  x"04",  x"04",  x"34",  x"52",  x"51",  x"1c",  x"1b", -- 1A98
         x"04",  x"04",  x"04",  x"26",  x"38",  x"40",  x"41",  x"45", -- 1AA0
         x"41",  x"04",  x"04",  x"04",  x"26",  x"52",  x"51",  x"04", -- 1AA8
         x"04",  x"04",  x"04",  x"26",  x"54",  x"53",  x"04",  x"04", -- 1AB0
         x"45",  x"41",  x"36",  x"35",  x"54",  x"53",  x"bf",  x"45", -- 1AB8
         x"04",  x"04",  x"04",  x"45",  x"15",  x"15",  x"14",  x"3d", -- 1AC0
         x"48",  x"04",  x"04",  x"04",  x"34",  x"54",  x"53",  x"42", -- 1AC8
         x"41",  x"42",  x"41",  x"45",  x"52",  x"51",  x"bf",  x"45", -- 1AD0
         x"15",  x"15",  x"37",  x"04",  x"52",  x"51",  x"be",  x"b2", -- 1AD8
         x"04",  x"04",  x"04",  x"47",  x"2f",  x"39",  x"43",  x"04", -- 1AE0
         x"04",  x"04",  x"04",  x"36",  x"35",  x"52",  x"51",  x"2c", -- 1AE8
         x"19",  x"15",  x"15",  x"58",  x"54",  x"53",  x"be",  x"b2", -- 1AF0
         x"5c",  x"3d",  x"43",  x"34",  x"54",  x"53",  x"27",  x"45", -- 1AF8
         x"45",  x"42",  x"41",  x"36",  x"35",  x"51",  x"45",  x"42", -- 1B00
         x"42",  x"41",  x"04",  x"45",  x"41",  x"54",  x"53",  x"18", -- 1B08
         x"15",  x"15",  x"15",  x"58",  x"52",  x"51",  x"45",  x"40", -- 1B10
         x"15",  x"41",  x"42",  x"40",  x"42",  x"40",  x"41",  x"47", -- 1B18
         x"15",  x"15",  x"15",  x"40",  x"41",  x"38",  x"15",  x"15", -- 1B20
         x"15",  x"14",  x"42",  x"15",  x"15",  x"40",  x"40",  x"42", -- 1B28
         x"17",  x"3d",  x"48",  x"47",  x"40",  x"40",  x"16",  x"15", -- 1B30
         x"19",  x"5d",  x"15",  x"15",  x"15",  x"15",  x"14",  x"41", -- 1B38
         x"15",  x"15",  x"15",  x"15",  x"18",  x"15",  x"15",  x"15", -- 1B40
         x"15",  x"13",  x"15",  x"15",  x"5c",  x"14",  x"15",  x"15", -- 1B48
         x"48",  x"04",  x"04",  x"45",  x"39",  x"15",  x"18",  x"19", -- 1B50
         x"15",  x"15",  x"5d",  x"19",  x"5d",  x"14",  x"15",  x"15", -- 1B58
         x"15",  x"15",  x"15",  x"15",  x"15",  x"16",  x"5c",  x"5c", -- 1B60
         x"14",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15",  x"18", -- 1B68
         x"42",  x"42",  x"41",  x"15",  x"40",  x"15",  x"18",  x"15", -- 1B70
         x"15",  x"15",  x"15",  x"15",  x"15",  x"13",  x"15",  x"15", -- 1B78
         x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 1B80
         x"15",  x"15",  x"14",  x"15",  x"15",  x"15",  x"15",  x"15", -- 1B88
         x"16",  x"15",  x"15",  x"5d",  x"15",  x"15",  x"19",  x"15", -- 1B90
         x"15",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15", -- 1B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1BC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1BC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1BD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc", -- 1BD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1BE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1BE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1BF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd", -- 1BF8
         x"00",  x"aa",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C10
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1C28
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C38
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1C48
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C50
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1C68
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C78
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C80
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C88
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C90
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C98
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CA0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CA8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CB0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CB8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CC0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CC8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CD0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CD8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CE0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CE8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CF0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CF8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D00
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D08
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D10
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D18
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D20
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D28
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D30
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D38
         x"15",  x"15",  x"5d",  x"21",  x"39",  x"15",  x"15",  x"15", -- 1D40
         x"13",  x"15",  x"14",  x"15",  x"15",  x"15",  x"15",  x"13", -- 1D48
         x"15",  x"15",  x"13",  x"15",  x"15",  x"2f",  x"22",  x"20", -- 1D50
         x"18",  x"15",  x"15",  x"13",  x"21",  x"22",  x"22",  x"20", -- 1D58
         x"15",  x"15",  x"14",  x"58",  x"52",  x"39",  x"5c",  x"14", -- 1D60
         x"16",  x"14",  x"16",  x"15",  x"15",  x"5c",  x"14",  x"15", -- 1D68
         x"4d",  x"14",  x"15",  x"15",  x"14",  x"54",  x"53",  x"2c", -- 1D70
         x"15",  x"16",  x"14",  x"15",  x"58",  x"54",  x"53",  x"2c", -- 1D78
         x"12",  x"11",  x"12",  x"4d",  x"54",  x"53",  x"2c",  x"4d", -- 1D80
         x"15",  x"15",  x"14",  x"18",  x"14",  x"15",  x"15",  x"11", -- 1D88
         x"0b",  x"10",  x"4d",  x"14",  x"58",  x"52",  x"51",  x"16", -- 1D90
         x"5c",  x"14",  x"17",  x"15",  x"58",  x"52",  x"51",  x"2c", -- 1D98
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"11",  x"0b", -- 1DA0
         x"12",  x"11",  x"12",  x"4d",  x"11",  x"10",  x"11",  x"0b", -- 1DA8
         x"0b",  x"0b",  x"0b",  x"12",  x"11",  x"54",  x"53",  x"11", -- 1DB0
         x"12",  x"4d",  x"11",  x"12",  x"4d",  x"54",  x"53",  x"11", -- 1DB8
         x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b", -- 1DC0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1DC8
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23", -- 1DD0
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23", -- 1DD8
         x"0b",  x"0b",  x"0b",  x"0b",  x"52",  x"51",  x"0b",  x"0b", -- 1DE0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1DE8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"0b", -- 1DF0
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"0b", -- 1DF8
         x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"38",  x"29",  x"30", -- 1E00
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1E08
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23", -- 1E10
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"52",  x"51",  x"23", -- 1E18
         x"0b",  x"0b",  x"0b",  x"10",  x"52",  x"39",  x"2c",  x"28", -- 1E20
         x"0b",  x"0b",  x"0b",  x"2a",  x"c1",  x"0b",  x"0b",  x"0b", -- 1E28
         x"c0",  x"c1",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"0b", -- 1E30
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"38",  x"29", -- 1E38
         x"c1",  x"0b",  x"2a",  x"c1",  x"54",  x"53",  x"28",  x"2a", -- 1E40
         x"c1",  x"c0",  x"1b",  x"04",  x"04",  x"1b",  x"1f",  x"c0", -- 1E48
         x"04",  x"04",  x"1f",  x"2a",  x"c1",  x"52",  x"51",  x"23", -- 1E50
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"39",  x"4d", -- 1E58
         x"04",  x"1b",  x"04",  x"26",  x"52",  x"51",  x"1b",  x"04", -- 1E60
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"1c",  x"04", -- 1E68
         x"04",  x"04",  x"1c",  x"04",  x"04",  x"54",  x"53",  x"c1", -- 1E70
         x"0b",  x"2a",  x"c1",  x"c0",  x"c1",  x"54",  x"53",  x"23", -- 1E78
         x"04",  x"04",  x"45",  x"42",  x"54",  x"53",  x"27",  x"04", -- 1E80
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1E88
         x"04",  x"45",  x"42",  x"41",  x"34",  x"52",  x"51",  x"27", -- 1E90
         x"1b",  x"04",  x"04",  x"04",  x"04",  x"52",  x"51",  x"1b", -- 1E98
         x"04",  x"04",  x"47",  x"58",  x"52",  x"51",  x"42",  x"41", -- 1EA0
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1EA8
         x"04",  x"47",  x"18",  x"5d",  x"40",  x"54",  x"53",  x"04", -- 1EB0
         x"04",  x"04",  x"04",  x"04",  x"34",  x"54",  x"53",  x"04", -- 1EB8
         x"04",  x"04",  x"04",  x"47",  x"54",  x"38",  x"15",  x"43", -- 1EC0
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1EC8
         x"04",  x"04",  x"47",  x"3d",  x"48",  x"52",  x"51",  x"bf", -- 1ED0
         x"04",  x"04",  x"04",  x"36",  x"35",  x"52",  x"51",  x"27", -- 1ED8
         x"04",  x"04",  x"04",  x"26",  x"52",  x"39",  x"43",  x"04", -- 1EE0
         x"04",  x"04",  x"45",  x"42",  x"41",  x"04",  x"04",  x"04", -- 1EE8
         x"04",  x"04",  x"04",  x"04",  x"34",  x"54",  x"53",  x"be", -- 1EF0
         x"bf",  x"04",  x"04",  x"04",  x"26",  x"54",  x"53",  x"27", -- 1EF8
         x"04",  x"04",  x"04",  x"34",  x"54",  x"53",  x"bf",  x"45", -- 1F00
         x"42",  x"42",  x"16",  x"5c",  x"14",  x"42",  x"41",  x"04", -- 1F08
         x"04",  x"45",  x"41",  x"36",  x"35",  x"52",  x"51",  x"45", -- 1F10
         x"19",  x"42",  x"42",  x"41",  x"45",  x"38",  x"40",  x"41", -- 1F18
         x"45",  x"41",  x"34",  x"35",  x"be",  x"38",  x"40",  x"5c", -- 1F20
         x"15",  x"15",  x"14",  x"15",  x"15",  x"15",  x"15",  x"41", -- 1F28
         x"45",  x"15",  x"15",  x"37",  x"45",  x"38",  x"40",  x"19", -- 1F30
         x"15",  x"15",  x"15",  x"19",  x"58",  x"39",  x"15",  x"15", -- 1F38
         x"5c",  x"14",  x"40",  x"42",  x"42",  x"16",  x"14",  x"15", -- 1F40
         x"17",  x"14",  x"5d",  x"19",  x"5d",  x"15",  x"15",  x"15", -- 1F48
         x"13",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"16", -- 1F50
         x"15",  x"15",  x"19",  x"15",  x"15",  x"40",  x"15",  x"15", -- 1F58
         x"15",  x"15",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15", -- 1F60
         x"15",  x"15",  x"15",  x"15",  x"15",  x"13",  x"15",  x"43", -- 1F68
         x"47",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 1F70
         x"17",  x"5c",  x"17",  x"15",  x"15",  x"15",  x"15",  x"15", -- 1F78
         x"15",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15", -- 1F80
         x"15",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"41", -- 1F88
         x"45",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 1F90
         x"15",  x"14",  x"15",  x"16",  x"15",  x"15",  x"15",  x"15", -- 1F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1FC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1FC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1FD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3", -- 1FD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1FE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1FE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1FF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
