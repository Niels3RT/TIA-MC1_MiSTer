library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_g4 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_g4;

architecture rtl of rom_g4 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"00",  x"ab",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0000
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0010
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0028
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0038
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0048
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0050
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0068
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0078
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0080
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0088
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0090
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0098
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 00A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 00A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 00B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 00B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 00C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 00C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 00D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 00D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 00E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 00E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 00F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 00F8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"67",  x"66", -- 0100
         x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03", -- 0108
         x"03",  x"03",  x"03",  x"03",  x"6c",  x"6b",  x"56",  x"56", -- 0110
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0118
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"6f",  x"6d", -- 0120
         x"68",  x"68",  x"68",  x"68",  x"68",  x"68",  x"68",  x"68", -- 0128
         x"68",  x"68",  x"68",  x"68",  x"6d",  x"6a",  x"55",  x"55", -- 0130
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0138
         x"15",  x"15",  x"15",  x"21",  x"22",  x"22",  x"20",  x"15", -- 0140
         x"15",  x"13",  x"15",  x"15",  x"5c",  x"2f",  x"22",  x"20", -- 0148
         x"17",  x"15",  x"15",  x"15",  x"5d",  x"15",  x"15",  x"21", -- 0150
         x"22",  x"22",  x"20",  x"15",  x"15",  x"17",  x"15",  x"15", -- 0158
         x"15",  x"15",  x"15",  x"14",  x"52",  x"51",  x"2c",  x"5c", -- 0160
         x"14",  x"16",  x"4d",  x"14",  x"15",  x"54",  x"53",  x"15", -- 0168
         x"14",  x"16",  x"5c",  x"14",  x"15",  x"15",  x"14",  x"16", -- 0170
         x"54",  x"53",  x"2c",  x"15",  x"15",  x"15",  x"16",  x"15", -- 0178
         x"12",  x"4d",  x"14",  x"58",  x"54",  x"53",  x"11",  x"12", -- 0180
         x"4d",  x"11",  x"0b",  x"10",  x"4d",  x"52",  x"51",  x"11", -- 0188
         x"12",  x"15",  x"15",  x"15",  x"15",  x"11",  x"12",  x"4d", -- 0190
         x"52",  x"51",  x"15",  x"15",  x"15",  x"4d",  x"11",  x"12", -- 0198
         x"0b",  x"0b",  x"12",  x"4d",  x"52",  x"51",  x"0b",  x"0b", -- 01A0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"38",  x"30", -- 01A8
         x"10",  x"11",  x"12",  x"4d",  x"11",  x"0b",  x"0b",  x"69", -- 01B0
         x"54",  x"53",  x"12",  x"4d",  x"11",  x"0b",  x"0b",  x"10", -- 01B8
         x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b", -- 01C0
         x"0b",  x"0b",  x"0b",  x"0b",  x"10",  x"52",  x"39",  x"28", -- 01C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69", -- 01D0
         x"52",  x"51",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 01D8
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b", -- 01E0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"c5",  x"c5",  x"0b", -- 01E8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 01F0
         x"54",  x"53",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 01F8
         x"0b",  x"0b",  x"0b",  x"10",  x"54",  x"38",  x"29",  x"30", -- 0200
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0208
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69", -- 0210
         x"52",  x"51",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0218
         x"0b",  x"0b",  x"0b",  x"0b",  x"52",  x"39",  x"15",  x"28", -- 0220
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0228
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69", -- 0230
         x"54",  x"53",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0238
         x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"28",  x"0b", -- 0240
         x"c0",  x"c1",  x"c0",  x"c1",  x"0b",  x"c0",  x"c1",  x"0b", -- 0248
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0250
         x"52",  x"51",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0258
         x"c0",  x"c1",  x"0b",  x"69",  x"52",  x"51",  x"1f",  x"c0", -- 0260
         x"04",  x"04",  x"04",  x"04",  x"1b",  x"04",  x"04",  x"1f", -- 0268
         x"2a",  x"1f",  x"c0",  x"c1",  x"0b",  x"2a",  x"c1",  x"69", -- 0270
         x"54",  x"53",  x"c1",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0278
         x"04",  x"04",  x"1b",  x"1b",  x"54",  x"53",  x"1c",  x"04", -- 0280
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"1c", -- 0288
         x"04",  x"1c",  x"04",  x"04",  x"1b",  x"04",  x"04",  x"1b", -- 0290
         x"38",  x"40",  x"41",  x"c1",  x"0b",  x"2a",  x"c1",  x"c0", -- 0298
         x"04",  x"04",  x"04",  x"26",  x"52",  x"51",  x"bf",  x"04", -- 02A0
         x"c4",  x"c2",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 02A8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"45", -- 02B0
         x"15",  x"15",  x"15",  x"41",  x"1b",  x"04",  x"04",  x"04", -- 02B8
         x"04",  x"04",  x"04",  x"04",  x"54",  x"53",  x"be",  x"04", -- 02C0
         x"04",  x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"04", -- 02C8
         x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"45",  x"16", -- 02D0
         x"2f",  x"39",  x"3d",  x"43",  x"04",  x"04",  x"04",  x"04", -- 02D8
         x"04",  x"c4",  x"c2",  x"34",  x"52",  x"51",  x"04",  x"04", -- 02E0
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 02E8
         x"c4",  x"c2",  x"04",  x"04",  x"04",  x"04",  x"47",  x"3d", -- 02F0
         x"54",  x"38",  x"41",  x"04",  x"04",  x"45",  x"41",  x"04", -- 02F8
         x"41",  x"04",  x"36",  x"35",  x"54",  x"53",  x"bf",  x"45", -- 0300
         x"42",  x"41",  x"45",  x"42",  x"42",  x"41",  x"04",  x"04", -- 0308
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"34", -- 0310
         x"52",  x"39",  x"43",  x"45",  x"42",  x"15",  x"15",  x"41", -- 0318
         x"15",  x"41",  x"04",  x"34",  x"52",  x"51",  x"be",  x"b2", -- 0320
         x"19",  x"5d",  x"15",  x"15",  x"15",  x"15",  x"42",  x"41", -- 0328
         x"04",  x"04",  x"04",  x"04",  x"45",  x"41",  x"36",  x"35", -- 0330
         x"be",  x"38",  x"42",  x"5d",  x"19",  x"15",  x"15",  x"15", -- 0338
         x"5d",  x"19",  x"42",  x"40",  x"40",  x"40",  x"41",  x"40", -- 0340
         x"15",  x"15",  x"5d",  x"19",  x"5d",  x"15",  x"15",  x"48", -- 0348
         x"04",  x"45",  x"41",  x"45",  x"15",  x"15",  x"40",  x"41", -- 0350
         x"45",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15", -- 0358
         x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0360
         x"15",  x"15",  x"14",  x"5c",  x"14",  x"19",  x"5d",  x"41", -- 0368
         x"45",  x"15",  x"15",  x"5d",  x"15",  x"15",  x"15",  x"15", -- 0370
         x"5d",  x"15",  x"15",  x"15",  x"19",  x"5d",  x"15",  x"15", -- 0378
         x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0380
         x"15",  x"14",  x"14",  x"15",  x"15",  x"15",  x"13",  x"14", -- 0388
         x"16",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15",  x"15", -- 0390
         x"14",  x"15",  x"15",  x"19",  x"15",  x"15",  x"5d",  x"15", -- 0398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03B8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 03C0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 03C8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 03D0
         x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3", -- 03D8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 03E0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 03E8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 03F0
         x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0", -- 03F8
         x"00",  x"ac",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0400
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0408
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0410
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0418
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0420
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0428
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0430
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0438
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0440
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0448
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0450
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0458
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0460
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0468
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0470
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0478
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0480
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0488
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0490
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0498
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 04A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 04A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 04B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 04B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 04C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 04C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 04D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 04D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 04E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 04E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 04F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 04F8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0500
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0508
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0510
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0518
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0520
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0528
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0530
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0538
         x"22",  x"20",  x"18",  x"15",  x"15",  x"15",  x"13",  x"15", -- 0540
         x"15",  x"15",  x"13",  x"15",  x"15",  x"15",  x"13",  x"15", -- 0548
         x"15",  x"13",  x"15",  x"17",  x"15",  x"17",  x"15",  x"17", -- 0550
         x"15",  x"15",  x"21",  x"22",  x"22",  x"20",  x"13",  x"15", -- 0558
         x"51",  x"2c",  x"15",  x"16",  x"5c",  x"14",  x"15",  x"15", -- 0560
         x"4d",  x"11",  x"12",  x"15",  x"15",  x"14",  x"16",  x"4d", -- 0568
         x"14",  x"15",  x"15",  x"15",  x"16",  x"4d",  x"16",  x"15", -- 0570
         x"16",  x"5c",  x"58",  x"52",  x"51",  x"14",  x"16",  x"13", -- 0578
         x"53",  x"15",  x"15",  x"14",  x"15",  x"16",  x"4d",  x"11", -- 0580
         x"0b",  x"0b",  x"0b",  x"10",  x"11",  x"12",  x"11",  x"0b", -- 0588
         x"10",  x"11",  x"12",  x"4d",  x"11",  x"0b",  x"10",  x"16", -- 0590
         x"5c",  x"14",  x"16",  x"54",  x"53",  x"12",  x"15",  x"15", -- 0598
         x"51",  x"10",  x"11",  x"12",  x"4d",  x"11",  x"0b",  x"0b", -- 05A0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 05A8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"10", -- 05B0
         x"11",  x"12",  x"11",  x"52",  x"51",  x"23",  x"12",  x"11", -- 05B8
         x"53",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 05C0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 05C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 05D0
         x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b",  x"0b", -- 05D8
         x"51",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 05E0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 05E8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 05F0
         x"0b",  x"0b",  x"0b",  x"52",  x"51",  x"0b",  x"0b",  x"0b", -- 05F8
         x"53",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0600
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0608
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0610
         x"0b",  x"0b",  x"69",  x"54",  x"53",  x"0b",  x"0b",  x"0b", -- 0618
         x"51",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0620
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0628
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0630
         x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b",  x"0b", -- 0638
         x"53",  x"30",  x"29",  x"29",  x"30",  x"33",  x"5e",  x"0b", -- 0640
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0648
         x"0b",  x"33",  x"5e",  x"0b",  x"0b",  x"0b",  x"24",  x"0b", -- 0650
         x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"23",  x"2a",  x"1f", -- 0658
         x"51",  x"2c",  x"16",  x"5c",  x"28",  x"25",  x"49",  x"5f", -- 0660
         x"5e",  x"1e",  x"1a",  x"9b",  x"1a",  x"0b",  x"2a",  x"1f", -- 0668
         x"0b",  x"2b",  x"49",  x"5f",  x"5e",  x"1e",  x"1d",  x"1e", -- 0670
         x"1a",  x"0b",  x"2a",  x"52",  x"51",  x"29",  x"41",  x"1c", -- 0678
         x"53",  x"15",  x"3d",  x"73",  x"49",  x"2e",  x"3b",  x"3c", -- 0680
         x"49",  x"2e",  x"03",  x"03",  x"4c",  x"1b",  x"04",  x"1c", -- 0688
         x"1b",  x"04",  x"3e",  x"01",  x"49",  x"2e",  x"03",  x"03", -- 0690
         x"4c",  x"1b",  x"26",  x"54",  x"38",  x"16",  x"14",  x"41", -- 0698
         x"51",  x"43",  x"04",  x"04",  x"5b",  x"5a",  x"4f",  x"4e", -- 06A0
         x"3e",  x"01",  x"2d",  x"4c",  x"04",  x"04",  x"04",  x"04", -- 06A8
         x"04",  x"04",  x"04",  x"3e",  x"01",  x"01",  x"2d",  x"4c", -- 06B0
         x"04",  x"04",  x"34",  x"52",  x"39",  x"15",  x"15",  x"14", -- 06B8
         x"53",  x"27",  x"45",  x"42",  x"41",  x"04",  x"04",  x"04", -- 06C0
         x"04",  x"3f",  x"4b",  x"04",  x"04",  x"04",  x"04",  x"04", -- 06C8
         x"04",  x"04",  x"04",  x"04",  x"3f",  x"4a",  x"4b",  x"45", -- 06D0
         x"41",  x"36",  x"35",  x"54",  x"53",  x"47",  x"48",  x"47", -- 06D8
         x"38",  x"42",  x"3a",  x"5d",  x"43",  x"04",  x"04",  x"04", -- 06E0
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 06E8
         x"04",  x"04",  x"45",  x"45",  x"41",  x"45",  x"42",  x"15", -- 06F0
         x"15",  x"37",  x"26",  x"52",  x"38",  x"41",  x"04",  x"04", -- 06F8
         x"15",  x"15",  x"15",  x"15",  x"15",  x"42",  x"42",  x"41", -- 0700
         x"45",  x"41",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0708
         x"04",  x"04",  x"47",  x"15",  x"14",  x"15",  x"15",  x"16", -- 0710
         x"3d",  x"43",  x"34",  x"54",  x"39",  x"43",  x"04",  x"04", -- 0718
         x"5d",  x"15",  x"15",  x"15",  x"19",  x"5d",  x"3d",  x"3d", -- 0720
         x"5c",  x"43",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0728
         x"04",  x"45",  x"42",  x"3a",  x"3a",  x"16",  x"19",  x"5d", -- 0730
         x"42",  x"42",  x"40",  x"40",  x"40",  x"41",  x"42",  x"41", -- 0738
         x"15",  x"41",  x"47",  x"14",  x"15",  x"15",  x"41",  x"45", -- 0740
         x"3a",  x"42",  x"41",  x"04",  x"04",  x"04",  x"04",  x"45", -- 0748
         x"42",  x"15",  x"15",  x"15",  x"15",  x"19",  x"15",  x"15", -- 0750
         x"5d",  x"19",  x"5d",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0758
         x"15",  x"15",  x"45",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0760
         x"15",  x"15",  x"43",  x"04",  x"04",  x"04",  x"04",  x"47", -- 0768
         x"15",  x"15",  x"15",  x"15",  x"19",  x"15",  x"15",  x"15", -- 0770
         x"15",  x"15",  x"15",  x"5d",  x"15",  x"15",  x"15",  x"15", -- 0778
         x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0780
         x"15",  x"15",  x"41",  x"04",  x"04",  x"04",  x"04",  x"45", -- 0788
         x"15",  x"15",  x"15",  x"3a",  x"15",  x"15",  x"15",  x"15", -- 0790
         x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15",  x"15", -- 0798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07B8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07C0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07C8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07D0
         x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07D8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07E0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07E8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07F0
         x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07F8
         x"00",  x"ad",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0810
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0828
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0838
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0848
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0850
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0868
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0878
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0880
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0888
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0890
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0898
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 08A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 08A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 08B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 08B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 08C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 08C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 08D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 08D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 08E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 08E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 08F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 08F8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0900
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0908
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0910
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0918
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0920
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0928
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0930
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0938
         x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"21",  x"22", -- 0940
         x"22",  x"20",  x"15",  x"15",  x"18",  x"15",  x"15",  x"15", -- 0948
         x"15",  x"17",  x"15",  x"18",  x"15",  x"15",  x"15",  x"15", -- 0950
         x"15",  x"15",  x"2f",  x"22",  x"20",  x"15",  x"15",  x"15", -- 0958
         x"16",  x"5c",  x"15",  x"15",  x"15",  x"14",  x"16",  x"52", -- 0960
         x"51",  x"15",  x"15",  x"15",  x"14",  x"16",  x"14",  x"16", -- 0968
         x"5c",  x"14",  x"16",  x"14",  x"16",  x"5c",  x"15",  x"15", -- 0970
         x"15",  x"14",  x"52",  x"51",  x"16",  x"5c",  x"5c",  x"14", -- 0978
         x"15",  x"15",  x"16",  x"4d",  x"11",  x"10",  x"58",  x"54", -- 0980
         x"53",  x"16",  x"4d",  x"14",  x"15",  x"14",  x"16",  x"4d", -- 0988
         x"15",  x"15",  x"4d",  x"11",  x"12",  x"15",  x"16",  x"5c", -- 0990
         x"14",  x"15",  x"54",  x"53",  x"2c",  x"14",  x"15",  x"15", -- 0998
         x"12",  x"4d",  x"11",  x"0b",  x"0b",  x"0b",  x"12",  x"52", -- 09A0
         x"51",  x"11",  x"0b",  x"12",  x"11",  x"12",  x"11",  x"0b", -- 09A8
         x"10",  x"11",  x"0b",  x"0b",  x"0b",  x"10",  x"4d",  x"4d", -- 09B0
         x"11",  x"12",  x"52",  x"51",  x"11",  x"12",  x"4d",  x"11", -- 09B8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54", -- 09C0
         x"53",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 09C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 09D0
         x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b",  x"0b",  x"0b", -- 09D8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52", -- 09E0
         x"51",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 09E8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 09F0
         x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b",  x"0b",  x"0b", -- 09F8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"54", -- 0A00
         x"53",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0A08
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0A10
         x"0b",  x"0b",  x"54",  x"53",  x"0b",  x"0b",  x"0b",  x"0b", -- 0A18
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52", -- 0A20
         x"51",  x"23",  x"0b",  x"33",  x"5e",  x"0b",  x"0b",  x"0b", -- 0A28
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0A30
         x"0b",  x"69",  x"52",  x"51",  x"c1",  x"0b",  x"0b",  x"0b", -- 0A38
         x"1d",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"54", -- 0A40
         x"53",  x"5f",  x"5e",  x"25",  x"49",  x"5f",  x"5e",  x"44", -- 0A48
         x"5e",  x"0b",  x"0b",  x"0b",  x"24",  x"0b",  x"0b",  x"0b", -- 0A50
         x"0b",  x"c0",  x"54",  x"53",  x"bf",  x"c1",  x"0b",  x"0b", -- 0A58
         x"03",  x"1d",  x"1e",  x"1a",  x"0b",  x"2a",  x"1b",  x"52", -- 0A60
         x"51",  x"5a",  x"49",  x"2e",  x"3b",  x"3c",  x"49",  x"01", -- 0A68
         x"49",  x"5f",  x"5e",  x"1e",  x"1d",  x"1e",  x"1a",  x"0b", -- 0A70
         x"2a",  x"26",  x"52",  x"51",  x"be",  x"bf",  x"1f",  x"0b", -- 0A78
         x"2e",  x"03",  x"03",  x"4c",  x"1b",  x"04",  x"26",  x"54", -- 0A80
         x"53",  x"27",  x"5b",  x"5a",  x"01",  x"2e",  x"3b",  x"3c", -- 0A88
         x"01",  x"01",  x"49",  x"2e",  x"03",  x"03",  x"4c",  x"1b", -- 0A90
         x"04",  x"36",  x"54",  x"53",  x"27",  x"04",  x"1c",  x"1b", -- 0A98
         x"01",  x"2d",  x"4c",  x"04",  x"04",  x"04",  x"36",  x"52", -- 0AA0
         x"51",  x"bf",  x"04",  x"04",  x"5b",  x"5a",  x"4f",  x"4e", -- 0AA8
         x"5b",  x"5a",  x"01",  x"01",  x"2d",  x"4c",  x"04",  x"04", -- 0AB0
         x"04",  x"26",  x"52",  x"51",  x"27",  x"04",  x"04",  x"04", -- 0AB8
         x"4a",  x"4b",  x"04",  x"c4",  x"c2",  x"04",  x"45",  x"54", -- 0AC0
         x"53",  x"be",  x"bf",  x"04",  x"04",  x"04",  x"04",  x"c4", -- 0AC8
         x"c2",  x"04",  x"3f",  x"4a",  x"4b",  x"04",  x"c4",  x"c2", -- 0AD0
         x"04",  x"34",  x"54",  x"53",  x"bf",  x"04",  x"04",  x"04", -- 0AD8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"47",  x"52", -- 0AE0
         x"38",  x"42",  x"40",  x"42",  x"42",  x"41",  x"04",  x"04", -- 0AE8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0AF0
         x"36",  x"35",  x"52",  x"51",  x"be",  x"04",  x"04",  x"04", -- 0AF8
         x"45",  x"42",  x"41",  x"04",  x"04",  x"04",  x"34",  x"54", -- 0B00
         x"39",  x"43",  x"47",  x"14",  x"16",  x"15",  x"41",  x"04", -- 0B08
         x"04",  x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"36", -- 0B10
         x"35",  x"26",  x"54",  x"53",  x"27",  x"04",  x"04",  x"04", -- 0B18
         x"17",  x"5c",  x"14",  x"42",  x"41",  x"36",  x"35",  x"38", -- 0B20
         x"40",  x"41",  x"45",  x"15",  x"15",  x"15",  x"14",  x"42", -- 0B28
         x"41",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B30
         x"04",  x"34",  x"52",  x"51",  x"04",  x"c4",  x"c3",  x"c2", -- 0B38
         x"15",  x"15",  x"15",  x"15",  x"14",  x"41",  x"45",  x"16", -- 0B40
         x"5c",  x"14",  x"5d",  x"19",  x"5d",  x"14",  x"15",  x"15", -- 0B48
         x"43",  x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"04", -- 0B50
         x"36",  x"35",  x"be",  x"53",  x"27",  x"04",  x"04",  x"04", -- 0B58
         x"15",  x"15",  x"5c",  x"14",  x"15",  x"15",  x"15",  x"15", -- 0B60
         x"15",  x"15",  x"15",  x"15",  x"15",  x"5d",  x"5c",  x"14", -- 0B68
         x"42",  x"41",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B70
         x"04",  x"04",  x"26",  x"52",  x"bf",  x"04",  x"04",  x"04", -- 0B78
         x"15",  x"14",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0B80
         x"15",  x"15",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15", -- 0B88
         x"15",  x"43",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B90
         x"04",  x"04",  x"34",  x"54",  x"be",  x"bf",  x"04",  x"04", -- 0B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0BC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0BC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc", -- 0BD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0BD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0BE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0BE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd", -- 0BF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0BF8
         x"00",  x"ae",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C10
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0C28
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C38
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0C48
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C50
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0C68
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C78
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C80
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C88
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C90
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C98
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 0CA0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 0CA8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 0CB0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 0CB8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 0CC0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 0CC8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 0CD0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 0CD8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 0CE0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 0CE8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 0CF0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 0CF8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0D00
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0D08
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0D10
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 0D18
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0D20
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0D28
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0D30
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 0D38
         x"15",  x"15",  x"15",  x"21",  x"22",  x"22",  x"20",  x"15", -- 0D40
         x"17",  x"15",  x"15",  x"15",  x"13",  x"15",  x"15",  x"13", -- 0D48
         x"15",  x"15",  x"2f",  x"22",  x"20",  x"15",  x"15",  x"18", -- 0D50
         x"15",  x"15",  x"15",  x"13",  x"21",  x"22",  x"22",  x"20", -- 0D58
         x"15",  x"15",  x"15",  x"58",  x"54",  x"53",  x"17",  x"15", -- 0D60
         x"15",  x"16",  x"5c",  x"14",  x"15",  x"15",  x"14",  x"15", -- 0D68
         x"5c",  x"14",  x"52",  x"51",  x"2c",  x"15",  x"15",  x"14", -- 0D70
         x"16",  x"5c",  x"14",  x"15",  x"58",  x"52",  x"51",  x"15", -- 0D78
         x"15",  x"4d",  x"4d",  x"14",  x"52",  x"51",  x"2c",  x"16", -- 0D80
         x"4d",  x"4d",  x"11",  x"12",  x"4d",  x"14",  x"15",  x"14", -- 0D88
         x"15",  x"58",  x"54",  x"53",  x"16",  x"5c",  x"14",  x"16", -- 0D90
         x"15",  x"15",  x"16",  x"4d",  x"14",  x"54",  x"53",  x"2c", -- 0D98
         x"11",  x"0b",  x"0b",  x"12",  x"54",  x"53",  x"4d",  x"11", -- 0DA0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"10",  x"11",  x"12", -- 0DA8
         x"4d",  x"11",  x"52",  x"51",  x"10",  x"4d",  x"4d",  x"11", -- 0DB0
         x"12",  x"4d",  x"11",  x"0b",  x"12",  x"52",  x"51",  x"4d", -- 0DB8
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b", -- 0DC0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0DC8
         x"0b",  x"0b",  x"54",  x"53",  x"23",  x"0b",  x"0b",  x"0b", -- 0DD0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"c5",  x"c5",  x"0b", -- 0DD8
         x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"23",  x"0b", -- 0DE0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0DE8
         x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b",  x"0b",  x"0b", -- 0DF0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0DF8
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b", -- 0E00
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0E08
         x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b",  x"0b",  x"0b", -- 0E10
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0E18
         x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"23",  x"0b", -- 0E20
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0E28
         x"0b",  x"0b",  x"52",  x"51",  x"23",  x"0b",  x"0b",  x"0b", -- 0E30
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 0E38
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b", -- 0E40
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"24",  x"0b",  x"0b", -- 0E48
         x"0b",  x"69",  x"54",  x"53",  x"0b",  x"0b",  x"0b",  x"0b", -- 0E50
         x"0b",  x"44",  x"5e",  x"0b",  x"0b",  x"24",  x"0b",  x"0b", -- 0E58
         x"1a",  x"9b",  x"1a",  x"69",  x"54",  x"53",  x"30",  x"44", -- 0E60
         x"5f",  x"5e",  x"44",  x"5e",  x"1e",  x"1d",  x"1e",  x"1a", -- 0E68
         x"9b",  x"1a",  x"52",  x"38",  x"29",  x"29",  x"30",  x"44", -- 0E70
         x"49",  x"01",  x"49",  x"5e",  x"1e",  x"1d",  x"1e",  x"1a", -- 0E78
         x"03",  x"03",  x"4c",  x"1b",  x"52",  x"51",  x"73",  x"01", -- 0E80
         x"3c",  x"49",  x"01",  x"49",  x"2e",  x"03",  x"03",  x"03", -- 0E88
         x"03",  x"4c",  x"54",  x"39",  x"5c",  x"5c",  x"73",  x"01", -- 0E90
         x"01",  x"01",  x"3c",  x"49",  x"2e",  x"03",  x"03",  x"4c", -- 0E98
         x"03",  x"4c",  x"04",  x"36",  x"54",  x"53",  x"bf",  x"3f", -- 0EA0
         x"4b",  x"3e",  x"01",  x"01",  x"01",  x"2e",  x"03",  x"03", -- 0EA8
         x"4c",  x"34",  x"52",  x"51",  x"15",  x"43",  x"04",  x"5b", -- 0EB0
         x"5a",  x"01",  x"2e",  x"3b",  x"01",  x"2d",  x"4c",  x"04", -- 0EB8
         x"4c",  x"04",  x"04",  x"26",  x"52",  x"51",  x"be",  x"04", -- 0EC0
         x"04",  x"04",  x"5b",  x"5a",  x"01",  x"01",  x"2d",  x"4c", -- 0EC8
         x"36",  x"35",  x"54",  x"53",  x"43",  x"04",  x"04",  x"04", -- 0ED0
         x"04",  x"5b",  x"5a",  x"4b",  x"3f",  x"4b",  x"04",  x"04", -- 0ED8
         x"04",  x"04",  x"04",  x"34",  x"54",  x"53",  x"27",  x"04", -- 0EE0
         x"04",  x"04",  x"04",  x"04",  x"3f",  x"4a",  x"4b",  x"04", -- 0EE8
         x"04",  x"26",  x"52",  x"51",  x"bf",  x"04",  x"04",  x"04", -- 0EF0
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0EF8
         x"42",  x"41",  x"36",  x"35",  x"52",  x"51",  x"bf",  x"04", -- 0F00
         x"04",  x"04",  x"04",  x"04",  x"45",  x"41",  x"04",  x"04", -- 0F08
         x"04",  x"34",  x"54",  x"53",  x"be",  x"bf",  x"04",  x"04", -- 0F10
         x"04",  x"04",  x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04", -- 0F18
         x"15",  x"15",  x"43",  x"26",  x"54",  x"53",  x"be",  x"bf", -- 0F20
         x"45",  x"41",  x"04",  x"45",  x"15",  x"14",  x"42",  x"41", -- 0F28
         x"34",  x"35",  x"52",  x"51",  x"45",  x"19",  x"42",  x"41", -- 0F30
         x"04",  x"04",  x"c4",  x"c2",  x"04",  x"04",  x"04",  x"04", -- 0F38
         x"5c",  x"16",  x"41",  x"45",  x"40",  x"40",  x"45",  x"40", -- 0F40
         x"15",  x"43",  x"45",  x"15",  x"15",  x"13",  x"15",  x"15", -- 0F48
         x"37",  x"45",  x"40",  x"40",  x"19",  x"15",  x"15",  x"14", -- 0F50
         x"42",  x"41",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0F58
         x"15",  x"5c",  x"14",  x"15",  x"15",  x"15",  x"5d",  x"15", -- 0F60
         x"15",  x"41",  x"47",  x"5c",  x"14",  x"15",  x"15",  x"15", -- 0F68
         x"19",  x"15",  x"15",  x"15",  x"16",  x"5c",  x"14",  x"15", -- 0F70
         x"15",  x"15",  x"41",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0F78
         x"14",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"16", -- 0F80
         x"15",  x"15",  x"45",  x"15",  x"15",  x"15",  x"15",  x"14", -- 0F88
         x"16",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15", -- 0F90
         x"15",  x"15",  x"43",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"fc", -- 0FB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0FC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0FC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3", -- 0FD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0FD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0FE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0FE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0", -- 0FF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0FF8
         x"00",  x"af",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1000
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1010
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1028
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1038
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1048
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1050
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1068
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1078
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1080
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1088
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1090
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1098
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 10A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 10A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 10B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 10B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 10C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 10C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 10D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 10D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 10E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 10E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 10F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 10F8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1100
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1108
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1110
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1118
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1120
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1128
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1130
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1138
         x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"13", -- 1140
         x"15",  x"15",  x"15",  x"15",  x"15",  x"2f",  x"22",  x"20", -- 1148
         x"17",  x"15",  x"15",  x"15",  x"13",  x"15",  x"5c",  x"13", -- 1150
         x"15",  x"17",  x"15",  x"15",  x"15",  x"15",  x"13",  x"15", -- 1158
         x"15",  x"15",  x"16",  x"14",  x"16",  x"5c",  x"14",  x"16", -- 1160
         x"5c",  x"5c",  x"14",  x"16",  x"58",  x"52",  x"51",  x"2c", -- 1168
         x"15",  x"16",  x"4d",  x"14",  x"16",  x"14",  x"15",  x"16", -- 1170
         x"5c",  x"14",  x"16",  x"5c",  x"5c",  x"14",  x"5c",  x"14", -- 1178
         x"12",  x"4d",  x"15",  x"15",  x"4d",  x"11",  x"12",  x"15", -- 1180
         x"15",  x"15",  x"15",  x"11",  x"12",  x"54",  x"53",  x"2c", -- 1188
         x"4d",  x"11",  x"0b",  x"12",  x"11",  x"12",  x"4d",  x"14", -- 1190
         x"15",  x"15",  x"58",  x"39",  x"5c",  x"14",  x"15",  x"15", -- 1198
         x"0b",  x"0b",  x"12",  x"11",  x"0b",  x"0b",  x"0b",  x"10", -- 11A0
         x"4d",  x"4d",  x"11",  x"0b",  x"69",  x"52",  x"51",  x"11", -- 11A8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"12", -- 11B0
         x"4d",  x"11",  x"12",  x"52",  x"39",  x"4d",  x"11",  x"12", -- 11B8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 11C0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"23", -- 11C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 11D0
         x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b",  x"0b", -- 11D8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 11E0
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b", -- 11E8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 11F0
         x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b",  x"0b", -- 11F8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1200
         x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"0b", -- 1208
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1210
         x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"23",  x"0b",  x"0b", -- 1218
         x"0b",  x"0b",  x"44",  x"5e",  x"0b",  x"0b",  x"0b",  x"24", -- 1220
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"52",  x"51",  x"23", -- 1228
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1230
         x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b",  x"0b", -- 1238
         x"5f",  x"49",  x"01",  x"49",  x"5f",  x"5e",  x"1e",  x"1d", -- 1240
         x"1e",  x"1a",  x"1e",  x"1a",  x"0b",  x"54",  x"53",  x"25", -- 1248
         x"5f",  x"5f",  x"5e",  x"44",  x"5e",  x"0b",  x"0b",  x"0b", -- 1250
         x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b",  x"0b", -- 1258
         x"01",  x"01",  x"01",  x"01",  x"01",  x"49",  x"2e",  x"03", -- 1260
         x"03",  x"03",  x"03",  x"4c",  x"1b",  x"52",  x"51",  x"bf", -- 1268
         x"3e",  x"01",  x"49",  x"01",  x"49",  x"5f",  x"5e",  x"1e", -- 1270
         x"1a",  x"9b",  x"1a",  x"52",  x"51",  x"1e",  x"1d",  x"1e", -- 1278
         x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"2d", -- 1280
         x"03",  x"03",  x"4c",  x"04",  x"34",  x"54",  x"53",  x"be", -- 1288
         x"bf",  x"3e",  x"01",  x"2e",  x"3c",  x"01",  x"49",  x"2e", -- 1290
         x"03",  x"03",  x"03",  x"54",  x"53",  x"01",  x"2e",  x"03", -- 1298
         x"3c",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"2d", -- 12A0
         x"03",  x"4c",  x"04",  x"36",  x"35",  x"52",  x"51",  x"27", -- 12A8
         x"be",  x"04",  x"3e",  x"01",  x"2e",  x"3b",  x"3c",  x"01", -- 12B0
         x"2e",  x"03",  x"03",  x"52",  x"51",  x"3e",  x"01",  x"2d", -- 12B8
         x"2e",  x"3b",  x"3c",  x"2e",  x"3c",  x"01",  x"01",  x"2d", -- 12C0
         x"4c",  x"04",  x"36",  x"35",  x"26",  x"54",  x"53",  x"27", -- 12C8
         x"04",  x"04",  x"04",  x"5b",  x"5a",  x"4f",  x"4e",  x"3e", -- 12D0
         x"01",  x"2d",  x"4c",  x"54",  x"53",  x"bf",  x"3f",  x"4b", -- 12D8
         x"5a",  x"4f",  x"4e",  x"3f",  x"4b",  x"3f",  x"4a",  x"4b", -- 12E0
         x"04",  x"04",  x"04",  x"04",  x"34",  x"52",  x"51",  x"04", -- 12E8
         x"c4",  x"c2",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 12F0
         x"3f",  x"4b",  x"26",  x"52",  x"51",  x"be",  x"bf",  x"04", -- 12F8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1300
         x"04",  x"04",  x"04",  x"04",  x"26",  x"54",  x"53",  x"27", -- 1308
         x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"04",  x"04", -- 1310
         x"04",  x"04",  x"34",  x"54",  x"53",  x"45",  x"40",  x"41", -- 1318
         x"04",  x"04",  x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04", -- 1320
         x"04",  x"04",  x"04",  x"04",  x"34",  x"52",  x"51",  x"bf", -- 1328
         x"04",  x"04",  x"04",  x"04",  x"04",  x"45",  x"42",  x"42", -- 1330
         x"41",  x"34",  x"35",  x"38",  x"40",  x"16",  x"15",  x"15", -- 1338
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1340
         x"c4",  x"c2",  x"04",  x"34",  x"35",  x"be",  x"53",  x"be", -- 1348
         x"bf",  x"04",  x"04",  x"04",  x"45",  x"15",  x"15",  x"15", -- 1350
         x"15",  x"37",  x"45",  x"15",  x"15",  x"15",  x"16",  x"15", -- 1358
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1360
         x"04",  x"04",  x"36",  x"35",  x"04",  x"26",  x"52",  x"04", -- 1368
         x"04",  x"04",  x"04",  x"04",  x"47",  x"3d",  x"15",  x"15", -- 1370
         x"15",  x"43",  x"47",  x"15",  x"15",  x"5c",  x"14",  x"15", -- 1378
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1380
         x"04",  x"04",  x"04",  x"04",  x"04",  x"34",  x"54",  x"27", -- 1388
         x"04",  x"04",  x"04",  x"04",  x"04",  x"45",  x"16",  x"15", -- 1390
         x"14",  x"41",  x"45",  x"16",  x"14",  x"15",  x"15",  x"15", -- 1398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13B8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 13C0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 13C8
         x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3", -- 13D0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 13D8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 13E0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 13E8
         x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0", -- 13F0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 13F8
         x"00",  x"b1",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1400
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1408
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1410
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1418
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1420
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1428
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1430
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1438
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1440
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1448
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1450
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1458
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1460
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1468
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1470
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1478
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1480
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1488
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1490
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1498
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14F8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1500
         x"67",  x"66",  x"03",  x"03",  x"03",  x"6c",  x"6b",  x"67", -- 1508
         x"66",  x"03",  x"03",  x"6c",  x"6b",  x"67",  x"66",  x"03", -- 1510
         x"03",  x"03",  x"6c",  x"6b",  x"56",  x"56",  x"56",  x"56", -- 1518
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1520
         x"6f",  x"6d",  x"68",  x"68",  x"68",  x"6d",  x"6a",  x"6f", -- 1528
         x"6d",  x"68",  x"68",  x"6d",  x"6a",  x"6f",  x"6d",  x"68", -- 1530
         x"68",  x"68",  x"6d",  x"6a",  x"55",  x"55",  x"55",  x"55", -- 1538
         x"15",  x"15",  x"13",  x"15",  x"16",  x"5c",  x"5c",  x"5c", -- 1540
         x"13",  x"16",  x"4d",  x"15",  x"15",  x"15",  x"15",  x"15", -- 1548
         x"15",  x"15",  x"15",  x"15",  x"16",  x"15",  x"15",  x"15", -- 1550
         x"15",  x"15",  x"14",  x"16",  x"15",  x"15",  x"5c",  x"14", -- 1558
         x"12",  x"14",  x"15",  x"15",  x"14",  x"15",  x"16",  x"14", -- 1560
         x"15",  x"11",  x"0b",  x"12",  x"11",  x"12",  x"15",  x"15", -- 1568
         x"5c",  x"14",  x"16",  x"4d",  x"14",  x"16",  x"4d",  x"5c", -- 1570
         x"5c",  x"14",  x"15",  x"58",  x"39",  x"14",  x"15",  x"15", -- 1578
         x"0b",  x"12",  x"4d",  x"11",  x"12",  x"4d",  x"4d",  x"4d", -- 1580
         x"11",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"12",  x"11", -- 1588
         x"12",  x"4d",  x"11",  x"0b",  x"12",  x"11",  x"0b",  x"12", -- 1590
         x"4d",  x"4d",  x"11",  x"12",  x"52",  x"39",  x"4d",  x"4d", -- 1598
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15A0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15A8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15B0
         x"0b",  x"0b",  x"0b",  x"69",  x"54",  x"53",  x"0b",  x"0b", -- 15B8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15C0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15D0
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"0b", -- 15D8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15E0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15E8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 15F0
         x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"0b",  x"0b", -- 15F8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1600
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1608
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1610
         x"0b",  x"0b",  x"0b",  x"69",  x"52",  x"51",  x"0b",  x"0b", -- 1618
         x"0b",  x"0b",  x"44",  x"5e",  x"0b",  x"0b",  x"44",  x"5e", -- 1620
         x"44",  x"5f",  x"5f",  x"5e",  x"0b",  x"44",  x"5e",  x"44", -- 1628
         x"5e",  x"44",  x"5e",  x"0b",  x"0b",  x"0b",  x"24",  x"0b", -- 1630
         x"0b",  x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"23",  x"0b", -- 1638
         x"5f",  x"5f",  x"01",  x"49",  x"5f",  x"5f",  x"01",  x"49", -- 1640
         x"2e",  x"3b",  x"3c",  x"49",  x"5f",  x"01",  x"49",  x"01", -- 1648
         x"49",  x"01",  x"49",  x"5f",  x"5e",  x"1e",  x"1d",  x"1e", -- 1650
         x"1d",  x"1e",  x"1a",  x"44",  x"52",  x"51",  x"1a",  x"9b", -- 1658
         x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01", -- 1660
         x"01",  x"2e",  x"03",  x"3b",  x"3c",  x"01",  x"01",  x"01", -- 1668
         x"01",  x"01",  x"01",  x"01",  x"49",  x"2d",  x"03",  x"03", -- 1670
         x"03",  x"03",  x"4c",  x"3e",  x"54",  x"53",  x"03",  x"03", -- 1678
         x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01",  x"01", -- 1680
         x"01",  x"01",  x"2e",  x"03",  x"03",  x"3b",  x"3c",  x"01", -- 1688
         x"2e",  x"3c",  x"01",  x"01",  x"01",  x"2d",  x"03",  x"03", -- 1690
         x"03",  x"4c",  x"04",  x"26",  x"52",  x"51",  x"03",  x"03", -- 1698
         x"01",  x"e5",  x"3c",  x"01",  x"01",  x"01",  x"01",  x"01", -- 16A0
         x"01",  x"01",  x"01",  x"2d",  x"03",  x"03",  x"4c",  x"3e", -- 16A8
         x"01",  x"2e",  x"3b",  x"3c",  x"01",  x"2e",  x"03",  x"03", -- 16B0
         x"4c",  x"04",  x"04",  x"26",  x"54",  x"53",  x"4f",  x"4e", -- 16B8
         x"3c",  x"01",  x"01",  x"e5",  x"3c",  x"01",  x"e5",  x"3c", -- 16C0
         x"01",  x"01",  x"01",  x"2d",  x"03",  x"4c",  x"04",  x"04", -- 16C8
         x"5b",  x"5a",  x"4f",  x"4e",  x"3e",  x"01",  x"2d",  x"4c", -- 16D0
         x"04",  x"04",  x"45",  x"42",  x"52",  x"51",  x"bf",  x"04", -- 16D8
         x"2e",  x"3b",  x"3c",  x"01",  x"2e",  x"3b",  x"3c",  x"2e", -- 16E0
         x"3c",  x"01",  x"01",  x"2d",  x"4c",  x"04",  x"04",  x"04", -- 16E8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"3f",  x"4b",  x"04", -- 16F0
         x"04",  x"04",  x"47",  x"3d",  x"54",  x"53",  x"be",  x"bf", -- 16F8
         x"5a",  x"4f",  x"4e",  x"5b",  x"5a",  x"4f",  x"4e",  x"3f", -- 1700
         x"4b",  x"3f",  x"4a",  x"4b",  x"04",  x"04",  x"c4",  x"c2", -- 1708
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1710
         x"04",  x"04",  x"04",  x"34",  x"52",  x"51",  x"45",  x"40", -- 1718
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1720
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1728
         x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"04",  x"45",  x"42", -- 1730
         x"42",  x"41",  x"34",  x"35",  x"38",  x"40",  x"16",  x"15", -- 1738
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1740
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1748
         x"04",  x"04",  x"04",  x"04",  x"04",  x"45",  x"15",  x"15", -- 1750
         x"15",  x"15",  x"37",  x"45",  x"15",  x"15",  x"15",  x"16", -- 1758
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1760
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1768
         x"04",  x"04",  x"04",  x"04",  x"04",  x"47",  x"3d",  x"15", -- 1770
         x"15",  x"15",  x"43",  x"47",  x"15",  x"15",  x"5c",  x"5c", -- 1778
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1780
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1788
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"45",  x"16", -- 1790
         x"15",  x"14",  x"41",  x"45",  x"16",  x"14",  x"15",  x"15", -- 1798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17B8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17C0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17C8
         x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17D0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17D8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17E0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17E8
         x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17F0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17F8
         x"00",  x"b0",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1810
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1828
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1838
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1848
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1850
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1868
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1878
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1880
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1888
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1890
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1898
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 18B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 18D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 18F8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1900
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1908
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1910
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1918
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1920
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1928
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1930
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1938
         x"5c",  x"15",  x"21",  x"22",  x"22",  x"20",  x"15",  x"15", -- 1940
         x"17",  x"15",  x"15",  x"13",  x"15",  x"15",  x"17",  x"15", -- 1948
         x"15",  x"15",  x"13",  x"21",  x"39",  x"15",  x"17",  x"15", -- 1950
         x"15",  x"15",  x"5c",  x"2f",  x"22",  x"20",  x"15",  x"15", -- 1958
         x"15",  x"16",  x"58",  x"54",  x"53",  x"2c",  x"15",  x"15", -- 1960
         x"15",  x"16",  x"15",  x"16",  x"4d",  x"5c",  x"14",  x"16", -- 1968
         x"4d",  x"14",  x"15",  x"58",  x"52",  x"39",  x"2c",  x"16", -- 1970
         x"5c",  x"14",  x"11",  x"52",  x"51",  x"15",  x"15",  x"15", -- 1978
         x"10",  x"11",  x"12",  x"52",  x"51",  x"10",  x"11",  x"12", -- 1980
         x"4d",  x"11",  x"12",  x"11",  x"0b",  x"12",  x"4d",  x"11", -- 1988
         x"0b",  x"12",  x"4d",  x"11",  x"54",  x"53",  x"12",  x"11", -- 1990
         x"12",  x"11",  x"0b",  x"c5",  x"c5",  x"12",  x"15",  x"15", -- 1998
         x"0b",  x"0b",  x"69",  x"54",  x"53",  x"23",  x"0b",  x"0b", -- 19A0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 19A8
         x"0b",  x"0b",  x"0b",  x"0b",  x"c5",  x"c5",  x"0b",  x"0b", -- 19B0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"12",  x"4d", -- 19B8
         x"0b",  x"0b",  x"0b",  x"52",  x"51",  x"0b",  x"0b",  x"0b", -- 19C0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 19C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 19D0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 19D8
         x"0b",  x"0b",  x"69",  x"54",  x"38",  x"30",  x"0b",  x"0b", -- 19E0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 19E8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 19F0
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 19F8
         x"0b",  x"0b",  x"10",  x"52",  x"39",  x"28",  x"0b",  x"0b", -- 1A00
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1A08
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1A10
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1A18
         x"0b",  x"0b",  x"0b",  x"54",  x"53",  x"0b",  x"0b",  x"0b", -- 1A20
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1A28
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1A30
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1A38
         x"24",  x"0b",  x"69",  x"52",  x"51",  x"23",  x"33",  x"5f", -- 1A40
         x"5e",  x"0b",  x"0b",  x"44",  x"5e",  x"0b",  x"33",  x"5e", -- 1A48
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"44",  x"5e",  x"9b", -- 1A50
         x"1a",  x"0b",  x"0b",  x"33",  x"5e",  x"0b",  x"0b",  x"0b", -- 1A58
         x"1d",  x"1e",  x"1a",  x"54",  x"53",  x"25",  x"01",  x"01", -- 1A60
         x"49",  x"5f",  x"5f",  x"01",  x"49",  x"5f",  x"01",  x"49", -- 1A68
         x"5f",  x"5e",  x"44",  x"5e",  x"44",  x"01",  x"49",  x"2e", -- 1A70
         x"03",  x"1a",  x"25",  x"01",  x"49",  x"5f",  x"5e",  x"0b", -- 1A78
         x"03",  x"03",  x"4c",  x"52",  x"51",  x"bf",  x"5b",  x"5a", -- 1A80
         x"01",  x"2e",  x"3b",  x"3c",  x"01",  x"01",  x"2e",  x"3b", -- 1A88
         x"3c",  x"49",  x"01",  x"49",  x"01",  x"01",  x"01",  x"01", -- 1A90
         x"2e",  x"03",  x"03",  x"3b",  x"3c",  x"01",  x"49",  x"5f", -- 1A98
         x"03",  x"4c",  x"26",  x"54",  x"53",  x"be",  x"42",  x"41", -- 1AA0
         x"5b",  x"5a",  x"4f",  x"4e",  x"3e",  x"01",  x"01",  x"2d", -- 1AA8
         x"03",  x"3b",  x"3c",  x"01",  x"01",  x"01",  x"01",  x"01", -- 1AB0
         x"01",  x"2e",  x"03",  x"03",  x"03",  x"3b",  x"3c",  x"01", -- 1AB8
         x"4c",  x"04",  x"36",  x"52",  x"51",  x"45",  x"15",  x"14", -- 1AC0
         x"42",  x"41",  x"04",  x"04",  x"04",  x"3e",  x"01",  x"2e", -- 1AC8
         x"03",  x"03",  x"4c",  x"5b",  x"5a",  x"01",  x"01",  x"01", -- 1AD0
         x"01",  x"01",  x"2d",  x"03",  x"03",  x"03",  x"4c",  x"3e", -- 1AD8
         x"04",  x"04",  x"26",  x"54",  x"38",  x"16",  x"14",  x"15", -- 1AE0
         x"3d",  x"43",  x"c4",  x"c3",  x"c2",  x"04",  x"3e",  x"01", -- 1AE8
         x"2d",  x"4c",  x"04",  x"04",  x"04",  x"3e",  x"2e",  x"3c", -- 1AF0
         x"01",  x"01",  x"2e",  x"03",  x"03",  x"4c",  x"04",  x"04", -- 1AF8
         x"04",  x"04",  x"34",  x"52",  x"39",  x"3d",  x"3d",  x"43", -- 1B00
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"3f", -- 1B08
         x"4b",  x"04",  x"04",  x"04",  x"04",  x"04",  x"3f",  x"4b", -- 1B10
         x"3e",  x"01",  x"01",  x"2d",  x"4c",  x"04",  x"04",  x"04", -- 1B18
         x"41",  x"34",  x"35",  x"54",  x"53",  x"27",  x"04",  x"04", -- 1B20
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B28
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B30
         x"04",  x"3f",  x"4a",  x"4b",  x"04",  x"04",  x"04",  x"04", -- 1B38
         x"15",  x"37",  x"41",  x"52",  x"51",  x"bf",  x"04",  x"04", -- 1B40
         x"45",  x"41",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B48
         x"c4",  x"c2",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B50
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B58
         x"15",  x"15",  x"58",  x"54",  x"53",  x"be",  x"bf",  x"45", -- 1B60
         x"15",  x"15",  x"41",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B68
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B70
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B78
         x"15",  x"15",  x"58",  x"52",  x"51",  x"45",  x"40",  x"15", -- 1B80
         x"15",  x"15",  x"14",  x"41",  x"04",  x"04",  x"04",  x"04", -- 1B88
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B90
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1BC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc", -- 1BC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1BD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1BD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1BE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd", -- 1BE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1BF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1BF8
         x"00",  x"9c",  x"a9",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C10
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1C28
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C38
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1C48
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C50
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1C68
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C78
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C80
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C88
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C90
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1C98
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CA0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CA8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CB0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 1CB8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CC0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CC8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CD0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 1CD8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CE0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CE8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CF0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 1CF8
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D00
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D08
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D10
         x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1D18
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D20
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D28
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D30
         x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1D38
         x"c6",  x"00",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1D40
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1D48
         x"12",  x"4d",  x"4d",  x"14",  x"15",  x"16",  x"21",  x"22", -- 1D50
         x"22",  x"20",  x"15",  x"15",  x"15",  x"15",  x"15",  x"15", -- 1D58
         x"c6",  x"00",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1D60
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1D68
         x"0b",  x"0b",  x"0b",  x"12",  x"4d",  x"14",  x"16",  x"52", -- 1D70
         x"51",  x"16",  x"5c",  x"15",  x"15",  x"15",  x"5c",  x"14", -- 1D78
         x"c6",  x"00",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1D80
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1D88
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"12",  x"4d",  x"54", -- 1D90
         x"53",  x"4d",  x"11",  x"10",  x"5c",  x"14",  x"15",  x"15", -- 1D98
         x"c6",  x"d5",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1DA0
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1DA8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"52", -- 1DB0
         x"51",  x"23",  x"0b",  x"0b",  x"12",  x"11",  x"12",  x"4d", -- 1DB8
         x"c6",  x"d3",  x"d2",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1DC0
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1DC8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54", -- 1DD0
         x"53",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1DD8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1DE0
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1DE8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"52", -- 1DF0
         x"51",  x"23",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1DF8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1E00
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1E08
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54", -- 1E10
         x"53",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1E18
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1E20
         x"c6",  x"c6",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1E28
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"52", -- 1E30
         x"38",  x"29",  x"30",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1E38
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1E40
         x"00",  x"07",  x"c6",  x"0b",  x"0b",  x"0b",  x"0b",  x"24", -- 1E48
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"69",  x"54", -- 1E50
         x"39",  x"15",  x"11",  x"0b",  x"0b",  x"0b",  x"0b",  x"0b", -- 1E58
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1E60
         x"00",  x"07",  x"c6",  x"49",  x"5f",  x"5e",  x"1e",  x"1d", -- 1E68
         x"1e",  x"1a",  x"9b",  x"1a",  x"0b",  x"2a",  x"c1",  x"52", -- 1E70
         x"51",  x"11",  x"0b",  x"0b",  x"0b",  x"44",  x"5f",  x"5e", -- 1E78
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1E80
         x"d5",  x"07",  x"c6",  x"3e",  x"01",  x"49",  x"2e",  x"03", -- 1E88
         x"03",  x"03",  x"03",  x"4c",  x"1b",  x"04",  x"34",  x"54", -- 1E90
         x"53",  x"1b",  x"c1",  x"c0",  x"1b",  x"5b",  x"5a",  x"49", -- 1E98
         x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c6",  x"c6", -- 1EA0
         x"d3",  x"d2",  x"c6",  x"04",  x"3e",  x"01",  x"01",  x"2e", -- 1EA8
         x"03",  x"03",  x"4c",  x"04",  x"04",  x"36",  x"35",  x"52", -- 1EB0
         x"51",  x"bf",  x"45",  x"42",  x"41",  x"04",  x"04",  x"5b", -- 1EB8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6", -- 1EC0
         x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"3e",  x"01",  x"01", -- 1EC8
         x"2d",  x"4c",  x"04",  x"04",  x"04",  x"45",  x"42",  x"54", -- 1ED0
         x"53",  x"be",  x"b2",  x"15",  x"15",  x"41",  x"04",  x"04", -- 1ED8
         x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"d1",  x"d0",  x"d0", -- 1EE0
         x"d0",  x"d0",  x"d0",  x"c9",  x"04",  x"04",  x"3f",  x"4a", -- 1EE8
         x"4b",  x"04",  x"45",  x"42",  x"42",  x"15",  x"58",  x"52", -- 1EF0
         x"51",  x"45",  x"15",  x"15",  x"15",  x"14",  x"42",  x"41", -- 1EF8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6", -- 1F00
         x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"c4",  x"c2",  x"04", -- 1F08
         x"04",  x"04",  x"47",  x"15",  x"15",  x"15",  x"15",  x"40", -- 1F10
         x"40",  x"15",  x"15",  x"15",  x"15",  x"13",  x"15",  x"15", -- 1F18
         x"04",  x"c4",  x"c2",  x"04",  x"04",  x"c6",  x"c6",  x"c6", -- 1F20
         x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"04",  x"04", -- 1F28
         x"45",  x"41",  x"45",  x"16",  x"15",  x"15",  x"15",  x"5c", -- 1F30
         x"14",  x"16",  x"5c",  x"5c",  x"14",  x"15",  x"15",  x"14", -- 1F38
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6", -- 1F40
         x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"04",  x"45", -- 1F48
         x"15",  x"15",  x"15",  x"15",  x"16",  x"5c",  x"14",  x"15", -- 1F50
         x"15",  x"15",  x"15",  x"15",  x"15",  x"15",  x"43",  x"47", -- 1F58
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c8",  x"04",  x"c8", -- 1F60
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"04",  x"45",  x"15", -- 1F68
         x"15",  x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15", -- 1F70
         x"15",  x"15",  x"15",  x"15",  x"5c",  x"14",  x"41",  x"45", -- 1F78
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1F80
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"47",  x"15", -- 1F88
         x"15",  x"15",  x"15",  x"43",  x"47",  x"15",  x"15",  x"15", -- 1F90
         x"15",  x"15",  x"15",  x"14",  x"15",  x"15",  x"15",  x"15", -- 1F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1FC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3", -- 1FC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1FD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 1FD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1FE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0", -- 1FE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 1FF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
