library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_g5 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_g5;

architecture rtl of rom_g5 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"00",  x"a9",  x"a9",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0000
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0010
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0028
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0038
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0048
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0050
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0068
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0078
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0080
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0088
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0090
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0098
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 00A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 00A8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 00B0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 00B8
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 00C0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 00C8
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 00D0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 00D8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 00E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6", -- 00E8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 00F0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 00F8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"c6", -- 0100
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6", -- 0108
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"d7", -- 0110
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0118
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"c6", -- 0120
         x"cd",  x"cc",  x"c6",  x"c6",  x"cf",  x"c6",  x"c7",  x"c6", -- 0128
         x"cf",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"d7", -- 0130
         x"c6",  x"c6",  x"cd",  x"cc",  x"c6",  x"c6",  x"c6",  x"c6", -- 0138
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"c6", -- 0140
         x"cb",  x"ca",  x"c6",  x"c6",  x"ce",  x"c6",  x"c7",  x"c6", -- 0148
         x"ce",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"d7", -- 0150
         x"c6",  x"c6",  x"cb",  x"ca",  x"c6",  x"c6",  x"c6",  x"c6", -- 0158
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d6",  x"c6",  x"c6", -- 0160
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6", -- 0168
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d6",  x"d6", -- 0170
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0178
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0180
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6", -- 0188
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0190
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0198
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6", -- 01A8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01B0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01B8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01C0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6", -- 01C8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01D0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01D8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6", -- 01E8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01F0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 01F8
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 0200
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0208
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 0210
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0218
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"c6", -- 0220
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0228
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0230
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0238
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"c6", -- 0240
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0248
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0250
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0258
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"c6", -- 0260
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0268
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0270
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0278
         x"c7",  x"c6",  x"c6",  x"00",  x"07",  x"c6",  x"04",  x"c6", -- 0280
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0288
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0290
         x"d0",  x"c6",  x"07",  x"00",  x"c6",  x"c6",  x"c6",  x"c7", -- 0298
         x"c7",  x"c6",  x"c6",  x"00",  x"07",  x"c6",  x"04",  x"c6", -- 02A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 02A8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 02B0
         x"d0",  x"c6",  x"07",  x"00",  x"c6",  x"c6",  x"c6",  x"c7", -- 02B8
         x"c6",  x"c6",  x"c6",  x"d5",  x"07",  x"c6",  x"04",  x"c8", -- 02C0
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8", -- 02C8
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8", -- 02D0
         x"04",  x"c6",  x"07",  x"d4",  x"c6",  x"c6",  x"c6",  x"c6", -- 02D8
         x"c6",  x"c6",  x"c6",  x"d3",  x"d2",  x"c6",  x"04",  x"04", -- 02E0
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 02E8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 02F0
         x"04",  x"c6",  x"d3",  x"d2",  x"c6",  x"c6",  x"c6",  x"c6", -- 02F8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04", -- 0300
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"c4", -- 0308
         x"c2",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0310
         x"04",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0318
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04", -- 0320
         x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"04", -- 0328
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0330
         x"04",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0338
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04", -- 0340
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0348
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0350
         x"d1",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 0358
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"04", -- 0360
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0368
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0370
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0378
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0380
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0388
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0390
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03B8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 03C0
         x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3", -- 03C8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 03D0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 03D8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 03E0
         x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0", -- 03E8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 03F0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 03F8
         x"00",  x"aa",  x"a9",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0400
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0408
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0410
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0418
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0420
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0428
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0430
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0438
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0440
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0448
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0450
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0458
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0460
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0468
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0470
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0478
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0480
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0488
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0490
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0498
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 04A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 04A8
         x"c6",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 04B0
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 04B8
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 04C0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c6",  x"c6",  x"c6", -- 04C8
         x"c6",  x"00",  x"00",  x"00",  x"c7",  x"c7",  x"c7",  x"c7", -- 04D0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 04D8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 04E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 04E8
         x"c6",  x"00",  x"00",  x"00",  x"00",  x"00",  x"07",  x"c6", -- 04F0
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 04F8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0500
         x"c6",  x"d7",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 0508
         x"c6",  x"00",  x"00",  x"00",  x"00",  x"00",  x"07",  x"c6", -- 0510
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0518
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cd",  x"cc", -- 0520
         x"c6",  x"d7",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 0528
         x"c6",  x"00",  x"00",  x"00",  x"00",  x"00",  x"07",  x"c6", -- 0530
         x"d0",  x"cf",  x"c6",  x"cf",  x"c6",  x"cf",  x"c6",  x"c6", -- 0538
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cb",  x"ca", -- 0540
         x"c6",  x"d7",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 0548
         x"c6",  x"00",  x"00",  x"00",  x"00",  x"d5",  x"07",  x"c6", -- 0550
         x"d0",  x"ce",  x"c6",  x"ce",  x"c6",  x"ce",  x"c6",  x"c6", -- 0558
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0560
         x"c6",  x"d6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 0568
         x"c6",  x"00",  x"00",  x"00",  x"c6",  x"d3",  x"d2",  x"c6", -- 0570
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0578
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0580
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 0588
         x"c6",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0590
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0598
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 05A0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 05A8
         x"c7",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 05B0
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 05B8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 05C0
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"07",  x"00", -- 05C8
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 05D0
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 05D8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 05E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"07",  x"00", -- 05E8
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 05F0
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 05F8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0600
         x"cf",  x"c6",  x"c6",  x"cf",  x"d0",  x"c6",  x"07",  x"00", -- 0608
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0610
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0618
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0620
         x"ce",  x"c6",  x"c6",  x"ce",  x"d0",  x"c6",  x"07",  x"d4", -- 0628
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0630
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0638
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0640
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"d3",  x"d2", -- 0648
         x"c6",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0650
         x"d0",  x"33",  x"5f",  x"c6",  x"c6",  x"0b",  x"44",  x"c6", -- 0658
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0660
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6", -- 0668
         x"c6",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0670
         x"d0",  x"5b",  x"5a",  x"c6",  x"c6",  x"49",  x"01",  x"c6", -- 0678
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 0680
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0688
         x"c7",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0690
         x"d0",  x"d9",  x"d8",  x"c6",  x"c6",  x"db",  x"da",  x"c6", -- 0698
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 06A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"07",  x"00", -- 06A8
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 06B0
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 06B8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 06C0
         x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"07",  x"00", -- 06C8
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 06D0
         x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 06D8
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8", -- 06E0
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c6",  x"07",  x"00", -- 06E8
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 06F0
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8", -- 06F8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0700
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"07",  x"d4", -- 0708
         x"00",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0710
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0718
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c4",  x"c3",  x"c2", -- 0720
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"d3",  x"d2", -- 0728
         x"c6",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0730
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0738
         x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0740
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6", -- 0748
         x"c6",  x"00",  x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6", -- 0750
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0758
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0760
         x"04",  x"04",  x"04",  x"04",  x"d1",  x"d0",  x"d0",  x"d0", -- 0768
         x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 0770
         x"c9",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0778
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0780
         x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6",  x"c6", -- 0788
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0790
         x"c6",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 07B8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07C0
         x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07C8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07D0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 07D8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07E0
         x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07E8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07F0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 07F8
         x"00",  x"ab",  x"a9",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0810
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0828
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0838
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0848
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0850
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0868
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0878
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0880
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0888
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0890
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0898
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08A8
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08B0
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08B8
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 08C0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 08C8
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08D0
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 08D8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08E8
         x"c6",  x"c6",  x"d0",  x"07",  x"00",  x"c6",  x"c6",  x"c6", -- 08F0
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 08F8
         x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"c6",  x"c6", -- 0900
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0908
         x"c6",  x"c6",  x"d0",  x"07",  x"00",  x"c6",  x"c6",  x"c6", -- 0910
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0918
         x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"cd",  x"cc", -- 0920
         x"c6",  x"c6",  x"cf",  x"c6",  x"c6",  x"cf",  x"c6",  x"c6", -- 0928
         x"c6",  x"c6",  x"d0",  x"07",  x"d4",  x"c6",  x"c6",  x"c6", -- 0930
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0938
         x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"cb",  x"ca", -- 0940
         x"c6",  x"c6",  x"ce",  x"c6",  x"c6",  x"ce",  x"c6",  x"c6", -- 0948
         x"c6",  x"c6",  x"d0",  x"d3",  x"d2",  x"c6",  x"c6",  x"c6", -- 0950
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0958
         x"c6",  x"c6",  x"c6",  x"c6",  x"d6",  x"c6",  x"c6",  x"c6", -- 0960
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0968
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0970
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0978
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0980
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0988
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0990
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0998
         x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7",  x"c7", -- 09A0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 09A8
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 09B0
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 09B8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 09C0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 09C8
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"00", -- 09D0
         x"07",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 09D8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 09E0
         x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"c6",  x"c6",  x"c6", -- 09E8
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"00", -- 09F0
         x"07",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 09F8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cf", -- 0A00
         x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"cd",  x"cc",  x"c6", -- 0A08
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"d5", -- 0A10
         x"07",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A18
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"ce", -- 0A20
         x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"cb",  x"ca",  x"c6", -- 0A28
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"d3", -- 0A30
         x"d2",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A38
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A40
         x"c6",  x"c6",  x"c6",  x"d6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A48
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A50
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A58
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A60
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A68
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A70
         x"c6",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0A78
         x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7",  x"c7", -- 0A80
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0A88
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0A90
         x"c7",  x"c7",  x"d0",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 0A98
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0AA0
         x"c6",  x"47",  x"58",  x"52",  x"38",  x"c6",  x"c6",  x"c6", -- 0AA8
         x"c6",  x"c6",  x"d0",  x"07",  x"00",  x"00",  x"00",  x"00", -- 0AB0
         x"07",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0AB8
         x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0AC0
         x"c6",  x"04",  x"47",  x"54",  x"39",  x"c6",  x"c6",  x"c6", -- 0AC8
         x"c6",  x"c6",  x"d0",  x"07",  x"00",  x"00",  x"00",  x"00", -- 0AD0
         x"07",  x"c6",  x"d0",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0AD8
         x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04", -- 0AE0
         x"c8",  x"04",  x"26",  x"52",  x"51",  x"c8",  x"04",  x"c8", -- 0AE8
         x"04",  x"c8",  x"04",  x"07",  x"d4",  x"00",  x"00",  x"d5", -- 0AF0
         x"07",  x"c6",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8", -- 0AF8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B00
         x"04",  x"04",  x"34",  x"54",  x"53",  x"04",  x"04",  x"04", -- 0B08
         x"04",  x"04",  x"04",  x"d3",  x"d2",  x"c6",  x"c6",  x"d3", -- 0B10
         x"d2",  x"c6",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B18
         x"04",  x"04",  x"04",  x"04",  x"04",  x"45",  x"42",  x"42", -- 0B20
         x"41",  x"34",  x"35",  x"52",  x"51",  x"bf",  x"45",  x"42", -- 0B28
         x"42",  x"41",  x"04",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0B30
         x"c6",  x"c6",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B38
         x"04",  x"04",  x"04",  x"45",  x"42",  x"15",  x"15",  x"15", -- 0B40
         x"14",  x"37",  x"45",  x"40",  x"40",  x"40",  x"16",  x"5c", -- 0B48
         x"3d",  x"48",  x"d1",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 0B50
         x"d0",  x"d0",  x"c9",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B58
         x"04",  x"04",  x"45",  x"15",  x"15",  x"16",  x"5c",  x"14", -- 0B60
         x"15",  x"15",  x"5d",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0B68
         x"41",  x"04",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0B70
         x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B78
         x"04",  x"04",  x"47",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0B80
         x"15",  x"15",  x"14",  x"15",  x"15",  x"15",  x"15",  x"15", -- 0B88
         x"15",  x"41",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0B90
         x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"04",  x"04",  x"04", -- 0B98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0BB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc", -- 0BC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0BC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0BD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0BD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd", -- 0BE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0BE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0BF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0BF8
         x"00",  x"ac",  x"a9",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 0C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C10
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 0C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 0C28
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C38
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 0C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 0C48
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C50
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 0C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0C68
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0C78
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C80
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C88
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C90
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 0C98
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0CA0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0CA8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0CB0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0CB8
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0CC0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c6",  x"c6",  x"c6", -- 0CC8
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0CD0
         x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0CD8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0CE0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0CE8
         x"c6",  x"00",  x"07",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0CF0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0CF8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"c6", -- 0D00
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D08
         x"c6",  x"00",  x"07",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0D10
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D18
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"cd", -- 0D20
         x"cc",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D28
         x"cf",  x"d5",  x"07",  x"cf",  x"c6",  x"c7",  x"c6",  x"c6", -- 0D30
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cf",  x"c6",  x"c6", -- 0D38
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7",  x"c6",  x"cb", -- 0D40
         x"ca",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D48
         x"ce",  x"d3",  x"d2",  x"ce",  x"c6",  x"c7",  x"c6",  x"c6", -- 0D50
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"ce",  x"c6",  x"c6", -- 0D58
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d6",  x"c6",  x"c6", -- 0D60
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D68
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0D70
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D78
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D80
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D88
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0D90
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0D98
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 0DA0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c6",  x"c6",  x"c6", -- 0DA8
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0DB0
         x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0DB8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0DC0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0DC8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0DD0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0DD8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0DE0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0DE8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0DF0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0DF8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cf", -- 0E00
         x"c6",  x"cf",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"5e", -- 0E08
         x"1e",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0E10
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cf",  x"c6",  x"c7", -- 0E18
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"ce", -- 0E20
         x"c6",  x"ce",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"49", -- 0E28
         x"2e",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0E30
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"ce",  x"c6",  x"c7", -- 0E38
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0E40
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"db", -- 0E48
         x"da",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0E50
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0E58
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0E60
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0E68
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7",  x"c6",  x"c6", -- 0E70
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0E78
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 0E80
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0E88
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0E90
         x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 0E98
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0EA0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"3c",  x"01",  x"c6", -- 0EA8
         x"c6",  x"2e",  x"03",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0EB0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0EB8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0EC0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"2d",  x"3b",  x"c6", -- 0EC8
         x"c6",  x"01",  x"2d",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0ED0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0ED8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0EE0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"4a",  x"4b",  x"c6", -- 0EE8
         x"c6",  x"5a",  x"4f",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0EF0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0EF8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0F00
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d9",  x"d8",  x"c6", -- 0F08
         x"c6",  x"d9",  x"d8",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0F10
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0F18
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0F20
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0F28
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 0F30
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 0F38
         x"04",  x"c7",  x"d0",  x"c6",  x"d0",  x"c6",  x"d0",  x"c6", -- 0F40
         x"d0",  x"c6",  x"d0",  x"c6",  x"04",  x"c8",  x"04",  x"c8", -- 0F48
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c6",  x"d0",  x"c6", -- 0F50
         x"d0",  x"c6",  x"d0",  x"c6",  x"d0",  x"c6",  x"d0",  x"c7", -- 0F58
         x"04",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 0F60
         x"d0",  x"d0",  x"d0",  x"d0",  x"04",  x"04",  x"04",  x"04", -- 0F68
         x"04",  x"04",  x"04",  x"04",  x"04",  x"d0",  x"d0",  x"d0", -- 0F70
         x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 0F78
         x"04",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 0F80
         x"d0",  x"d0",  x"d0",  x"d0",  x"04",  x"04",  x"c4",  x"c3", -- 0F88
         x"c2",  x"04",  x"04",  x"04",  x"04",  x"d0",  x"d0",  x"d0", -- 0F90
         x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 0F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0FB8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3", -- 0FC0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0FC8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0FD0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 0FD8
         x"e1",  x"e0",  x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0", -- 0FE0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0FE8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0FF0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 0FF8
         x"00",  x"ad",  x"a9",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1000
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1010
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1028
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1038
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1048
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1050
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1068
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1078
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1080
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1088
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1090
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1098
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10A8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10B0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10B8
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 10C0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 10C8
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 10D0
         x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 10D8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10E8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10F0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 10F8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1100
         x"d7",  x"d7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1108
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1110
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d7", -- 1118
         x"c6",  x"c6",  x"cf",  x"c6",  x"c6",  x"cd",  x"cc",  x"c6", -- 1120
         x"d7",  x"d7",  x"c6",  x"cd",  x"cc",  x"c6",  x"c6",  x"c6", -- 1128
         x"c6",  x"c7",  x"c6",  x"cf",  x"c6",  x"c6",  x"c6",  x"c6", -- 1130
         x"c6",  x"c6",  x"c6",  x"c6",  x"cd",  x"cc",  x"c6",  x"d7", -- 1138
         x"c6",  x"c6",  x"ce",  x"c6",  x"c6",  x"cb",  x"ca",  x"c6", -- 1140
         x"d7",  x"d7",  x"c6",  x"cb",  x"ca",  x"c6",  x"c6",  x"c6", -- 1148
         x"c6",  x"c7",  x"c6",  x"ce",  x"c6",  x"c6",  x"c6",  x"c6", -- 1150
         x"c6",  x"c6",  x"c6",  x"c6",  x"cb",  x"ca",  x"c6",  x"d7", -- 1158
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1160
         x"d6",  x"d6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1168
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1170
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d6", -- 1178
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1180
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1188
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1190
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1198
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 11A0
         x"c7",  x"c7",  x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7", -- 11A8
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 11B0
         x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 11B8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 11C0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 11C8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 11D0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 11D8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 11E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 11E8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 11F0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 11F8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1200
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cf", -- 1208
         x"c6",  x"c6",  x"c6",  x"c6",  x"cf",  x"c6",  x"c6",  x"c6", -- 1210
         x"c6",  x"cf",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1218
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1220
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"ce", -- 1228
         x"c6",  x"c6",  x"c6",  x"c6",  x"ce",  x"c6",  x"c6",  x"c6", -- 1230
         x"c6",  x"ce",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1238
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1240
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1248
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1250
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1258
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7",  x"c7",  x"c7", -- 1260
         x"c7",  x"c7",  x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c7", -- 1268
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 1270
         x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7",  x"c7", -- 1278
         x"c6",  x"c7",  x"3b",  x"3c",  x"c6",  x"c6",  x"c6",  x"2e", -- 1280
         x"03",  x"c6",  x"c6",  x"c6",  x"d0",  x"d0",  x"c6",  x"c6", -- 1288
         x"c6",  x"d0",  x"d0",  x"c6",  x"c6",  x"c6",  x"d0",  x"d0", -- 1290
         x"c6",  x"c6",  x"c6",  x"d0",  x"d0",  x"c6",  x"c6",  x"c7", -- 1298
         x"c6",  x"c7",  x"2e",  x"03",  x"c6",  x"c6",  x"c6",  x"01", -- 12A0
         x"2d",  x"c6",  x"c6",  x"c6",  x"d0",  x"d0",  x"c6",  x"c6", -- 12A8
         x"c6",  x"d0",  x"d0",  x"c6",  x"c6",  x"c6",  x"d0",  x"d0", -- 12B0
         x"c6",  x"c6",  x"c6",  x"d0",  x"d0",  x"c6",  x"c6",  x"c7", -- 12B8
         x"c6",  x"c7",  x"4a",  x"4b",  x"c6",  x"c6",  x"c6",  x"5a", -- 12C0
         x"4f",  x"c6",  x"c6",  x"c6",  x"d0",  x"d0",  x"c6",  x"c6", -- 12C8
         x"c6",  x"d0",  x"d0",  x"c6",  x"c6",  x"c6",  x"d0",  x"d0", -- 12D0
         x"c6",  x"c6",  x"c6",  x"d0",  x"d0",  x"c6",  x"c6",  x"c7", -- 12D8
         x"c6",  x"c7",  x"d9",  x"d8",  x"c6",  x"c6",  x"c6",  x"d9", -- 12E0
         x"d8",  x"c6",  x"c6",  x"c6",  x"d3",  x"d2",  x"c6",  x"c6", -- 12E8
         x"c6",  x"d3",  x"d2",  x"c6",  x"c6",  x"c6",  x"d3",  x"d2", -- 12F0
         x"c6",  x"c6",  x"c6",  x"d3",  x"d2",  x"c6",  x"c6",  x"c7", -- 12F8
         x"c6",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1300
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1308
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1310
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1318
         x"c7",  x"c7",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1320
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1328
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1330
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c7", -- 1338
         x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8",  x"04",  x"c8", -- 1340
         x"04",  x"c8",  x"07",  x"c6",  x"d0",  x"c6",  x"d0",  x"c6", -- 1348
         x"d0",  x"c6",  x"d0",  x"c6",  x"d0",  x"c6",  x"d0",  x"c6", -- 1350
         x"d0",  x"c6",  x"07",  x"c6",  x"d0",  x"c6",  x"d0",  x"c6", -- 1358
         x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"04", -- 1360
         x"04",  x"04",  x"07",  x"d4",  x"d0",  x"d0",  x"d0",  x"d0", -- 1368
         x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 1370
         x"d0",  x"d5",  x"07",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 1378
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"c4",  x"c2", -- 1380
         x"04",  x"04",  x"d3",  x"d2",  x"d0",  x"d0",  x"d0",  x"d0", -- 1388
         x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 1390
         x"d0",  x"d3",  x"d2",  x"d0",  x"d0",  x"d0",  x"d0",  x"d0", -- 1398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 13B8
         x"e4",  x"e3",  x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3", -- 13C0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 13C8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 13D0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 13D8
         x"e1",  x"e0",  x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0", -- 13E0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 13E8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 13F0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 13F8
         x"00",  x"ae",  x"a9",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1400
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1408
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1410
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1418
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1420
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1428
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1430
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1438
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1440
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1448
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1450
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1458
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1460
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1468
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1470
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1478
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1480
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1488
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1490
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1498
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14A0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14A8
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14B0
         x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61",  x"61", -- 14B8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14C0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14C8
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14D0
         x"60",  x"59",  x"60",  x"59",  x"60",  x"59",  x"60",  x"59", -- 14D8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14E0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14E8
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14F0
         x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57",  x"57", -- 14F8
         x"56",  x"56",  x"56",  x"56",  x"67",  x"66",  x"03",  x"03", -- 1500
         x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03", -- 1508
         x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03", -- 1510
         x"03",  x"6c",  x"6b",  x"56",  x"56",  x"56",  x"56",  x"56", -- 1518
         x"55",  x"55",  x"55",  x"55",  x"6f",  x"6d",  x"68",  x"68", -- 1520
         x"68",  x"68",  x"68",  x"68",  x"68",  x"68",  x"68",  x"68", -- 1528
         x"68",  x"68",  x"68",  x"68",  x"68",  x"68",  x"68",  x"68", -- 1530
         x"68",  x"6d",  x"6a",  x"55",  x"55",  x"55",  x"55",  x"55", -- 1538
         x"15",  x"15",  x"15",  x"13",  x"15",  x"c6",  x"c6",  x"c6", -- 1540
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1548
         x"15",  x"5c",  x"14",  x"15",  x"c6",  x"c6",  x"c6",  x"16", -- 1550
         x"5c",  x"14",  x"15",  x"c6",  x"c6",  x"d0",  x"07",  x"00", -- 1558
         x"15",  x"15",  x"14",  x"16",  x"5c",  x"c6",  x"c6",  x"c6", -- 1560
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1568
         x"14",  x"15",  x"4d",  x"14",  x"c6",  x"c6",  x"c6",  x"15", -- 1570
         x"15",  x"16",  x"15",  x"c6",  x"c6",  x"d0",  x"07",  x"00", -- 1578
         x"5c",  x"14",  x"15",  x"11",  x"12",  x"c6",  x"c6",  x"c6", -- 1580
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1588
         x"12",  x"11",  x"0b",  x"12",  x"c6",  x"cf",  x"c6",  x"12", -- 1590
         x"4d",  x"11",  x"12",  x"c6",  x"c6",  x"d0",  x"07",  x"00", -- 1598
         x"12",  x"4d",  x"11",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6", -- 15A0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 15A8
         x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"ce",  x"c6",  x"0b", -- 15B0
         x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"d0",  x"07",  x"d4", -- 15B8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6", -- 15C0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 15C8
         x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6",  x"0b", -- 15D0
         x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"d0",  x"d3",  x"d2", -- 15D8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6", -- 15E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 15E8
         x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6",  x"0b", -- 15F0
         x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 15F8
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6", -- 1600
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1608
         x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6",  x"0b", -- 1610
         x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1618
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"07", -- 1620
         x"07",  x"07",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1628
         x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"c6",  x"0b", -- 1630
         x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1638
         x"0b",  x"0b",  x"0b",  x"0b",  x"0b",  x"c6",  x"c6",  x"07", -- 1640
         x"00",  x"00",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1648
         x"0b",  x"0b",  x"44",  x"5e",  x"c6",  x"c6",  x"c6",  x"5e", -- 1650
         x"0b",  x"0b",  x"44",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1658
         x"44",  x"5e",  x"0b",  x"0b",  x"44",  x"c6",  x"c6",  x"07", -- 1660
         x"00",  x"00",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1668
         x"5f",  x"49",  x"01",  x"49",  x"c6",  x"c6",  x"c6",  x"49", -- 1670
         x"5f",  x"49",  x"01",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1678
         x"01",  x"49",  x"5f",  x"49",  x"01",  x"c6",  x"c6",  x"07", -- 1680
         x"00",  x"00",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1688
         x"db",  x"01",  x"e5",  x"da",  x"c6",  x"c6",  x"c6",  x"db", -- 1690
         x"01",  x"01",  x"da",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 1698
         x"e5",  x"3c",  x"01",  x"e5",  x"3c",  x"c6",  x"c6",  x"07", -- 16A0
         x"d4",  x"d5",  x"07",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 16A8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 16B0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 16B8
         x"01",  x"2e",  x"3b",  x"3c",  x"2e",  x"c6",  x"c6",  x"d3", -- 16C0
         x"d2",  x"d3",  x"d2",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 16C8
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 16D0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"d0",  x"c6",  x"c6", -- 16D8
         x"5b",  x"5a",  x"4f",  x"4e",  x"3f",  x"c6",  x"c6",  x"c6", -- 16E0
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"c8",  x"04", -- 16E8
         x"c8",  x"5b",  x"c8",  x"4e",  x"c8",  x"04",  x"c8",  x"04", -- 16F0
         x"c8",  x"3e",  x"c8",  x"2d",  x"c8",  x"04",  x"c6",  x"c6", -- 16F8
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6", -- 1700
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"04", -- 1708
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1710
         x"04",  x"04",  x"3f",  x"4b",  x"04",  x"04",  x"c6",  x"c6", -- 1718
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6", -- 1720
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"c4", -- 1728
         x"c2",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1730
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6", -- 1738
         x"04",  x"04",  x"04",  x"c4",  x"c3",  x"c6",  x"c6",  x"c6", -- 1740
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04",  x"04", -- 1748
         x"04",  x"04",  x"c4",  x"c3",  x"c2",  x"04",  x"04",  x"04", -- 1750
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6", -- 1758
         x"04",  x"04",  x"04",  x"04",  x"d1",  x"d0",  x"d0",  x"d0", -- 1760
         x"d0",  x"d0",  x"d0",  x"d0",  x"d0",  x"c9",  x"04",  x"04", -- 1768
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1770
         x"04",  x"04",  x"04",  x"04",  x"04",  x"d1",  x"d0",  x"d0", -- 1778
         x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6",  x"c6", -- 1780
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"04",  x"04", -- 1788
         x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04",  x"04", -- 1790
         x"04",  x"04",  x"04",  x"04",  x"04",  x"c6",  x"c6",  x"c6", -- 1798
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 17B8
         x"e2",  x"dc",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17C0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17C8
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17D0
         x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3",  x"e4",  x"e3", -- 17D8
         x"de",  x"dd",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17E0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17E8
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17F0
         x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0",  x"e1",  x"e0", -- 17F8
         x"00",  x"9c",  x"9c",  x"a3",  x"a1",  x"a8",  x"a5",  x"b4", -- 1800
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1808
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1810
         x"00",  x"00",  x"9c",  x"9c",  x"a3",  x"9c",  x"9c",  x"00", -- 1818
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1820
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1828
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1830
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1838
         x"00",  x"9c",  x"9c",  x"a3",  x"b3",  x"b4",  x"ac",  x"9c", -- 1840
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1848
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1850
         x"00",  x"00",  x"b8",  x"50",  x"9e",  x"a1",  x"94",  x"00", -- 1858
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1860
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 1868
         x"df",  x"00",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1870
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1878
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1880
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1888
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1890
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1898
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 18F8
         x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1900
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1908
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1910
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"00",  x"00", -- 1918
         x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1920
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1928
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1930
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"00",  x"00", -- 1938
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1940
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1948
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1950
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1958
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1960
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1968
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1970
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1978
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1980
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1988
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1990
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1998
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 19A0
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 19A8
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 19B0
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 19B8
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 19C0
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 19C8
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 19D0
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 19D8
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 19E0
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 19E8
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 19F0
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 19F8
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1A00
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A08
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A10
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1A18
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1A20
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A28
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A30
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1A38
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1A40
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A48
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A50
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1A58
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1A60
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A68
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A70
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1A78
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1A80
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A88
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1A90
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1A98
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1AA0
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1AA8
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1AB0
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1AB8
         x"00",  x"00",  x"c6",  x"c6",  x"07",  x"07",  x"07",  x"07", -- 1AC0
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1AC8
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1AD0
         x"07",  x"07",  x"07",  x"07",  x"c6",  x"c6",  x"00",  x"00", -- 1AD8
         x"00",  x"00",  x"c6",  x"c6",  x"d3",  x"07",  x"07",  x"07", -- 1AE0
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1AE8
         x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07",  x"07", -- 1AF0
         x"07",  x"07",  x"07",  x"d2",  x"c6",  x"c6",  x"00",  x"00", -- 1AF8
         x"00",  x"00",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1B00
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"cd", -- 1B08
         x"cc",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6", -- 1B10
         x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"c6",  x"00",  x"00", -- 1B18
         x"00",  x"00",  x"c6",  x"00",  x"c6",  x"00",  x"c6",  x"00", -- 1B20
         x"c6",  x"00",  x"c6",  x"00",  x"c6",  x"00",  x"c6",  x"cb", -- 1B28
         x"ca",  x"c6",  x"00",  x"c6",  x"00",  x"c6",  x"00",  x"c6", -- 1B30
         x"00",  x"c6",  x"00",  x"c6",  x"00",  x"c6",  x"00",  x"00", -- 1B38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1B78
         x"00",  x"00",  x"79",  x"78",  x"7b",  x"7a",  x"81",  x"78", -- 1B80
         x"93",  x"92",  x"91",  x"90",  x"8b",  x"8a",  x"7b",  x"7a", -- 1B88
         x"00",  x"88",  x"9a",  x"99",  x"79",  x"78",  x"83",  x"82", -- 1B90
         x"81",  x"78",  x"7b",  x"7a",  x"79",  x"78",  x"00",  x"00", -- 1B98
         x"00",  x"00",  x"75",  x"74",  x"77",  x"76",  x"7d",  x"7c", -- 1BA0
         x"8f",  x"8e",  x"8d",  x"8c",  x"87",  x"84",  x"77",  x"76", -- 1BA8
         x"85",  x"84",  x"98",  x"97",  x"75",  x"74",  x"7f",  x"7e", -- 1BB0
         x"7d",  x"7c",  x"77",  x"76",  x"75",  x"74",  x"00",  x"00", -- 1BB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1BF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"65",  x"64",  x"65", -- 1C68
         x"64",  x"65",  x"64",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"63",  x"62",  x"63", -- 1C88
         x"62",  x"63",  x"62",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"71", -- 1CE0
         x"a5",  x"80",  x"9e",  x"a4",  x"6e",  x"a2",  x"00",  x"50", -- 1CE8
         x"a5",  x"94",  x"00",  x"50",  x"9e",  x"a5",  x"96",  x"9e", -- 1CF0
         x"95",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D30
         x"bc",  x"b3",  x"96",  x"9e",  x"70",  x"00",  x"00",  x"00", -- 1D38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"b3",  x"9c", -- 1D60
         x"9d",  x"9d",  x"9e",  x"ac",  x"9e",  x"50",  x"a5",  x"9d", -- 1D68
         x"00",  x"b4",  x"00",  x"b5",  x"6e",  x"9e",  x"a7",  x"b3", -- 1D70
         x"a5",  x"9f",  x"b3",  x"94",  x"a8",  x"00",  x"00",  x"00", -- 1D78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"bd",  x"bb",  x"00", -- 1D80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"bb", -- 1D90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"bc",  x"b8",  x"b3", -- 1DA0
         x"94",  x"a7",  x"6e",  x"a7",  x"b8",  x"a4",  x"9e",  x"a1", -- 1DA8
         x"a4",  x"00",  x"b8",  x"a5",  x"94",  x"9e",  x"96",  x"9c", -- 1DB0
         x"a8",  x"9c",  x"9e",  x"a1",  x"a4",  x"00",  x"00",  x"00", -- 1DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"bc",  x"ba", -- 1DF0
         x"b5",  x"a1",  x"a5",  x"a8",  x"a2",  x"00",  x"00",  x"00", -- 1DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E00
         x"00",  x"00",  x"00",  x"00",  x"bd",  x"00",  x"00",  x"00", -- 1E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"bd",  x"00",  x"00", -- 1E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E18
         x"00",  x"00",  x"00",  x"00",  x"b5",  x"a7",  x"b3",  x"6e", -- 1E20
         x"9c",  x"9d",  x"a5",  x"9d",  x"bc",  x"b8",  x"6e",  x"b5", -- 1E28
         x"a7",  x"b3",  x"95",  x"9c",  x"96",  x"bc",  x"b5",  x"a7", -- 1E30
         x"a5",  x"9f",  x"a6",  x"a1",  x"a4",  x"00",  x"00",  x"00", -- 1E38
         x"00",  x"00",  x"00",  x"00",  x"bd",  x"00",  x"00",  x"00", -- 1E40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E58
         x"00",  x"00",  x"00",  x"00",  x"bc",  x"a8",  x"a5",  x"ab", -- 1E60
         x"a5",  x"9d",  x"00",  x"b3",  x"00",  x"a8",  x"9e",  x"a1", -- 1E68
         x"9e",  x"a4",  x"94",  x"00",  x"b8",  x"6e",  x"b5",  x"a7", -- 1E70
         x"a5",  x"9f",  x"b3",  x"94",  x"a8",  x"00",  x"00",  x"00", -- 1E78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E98
         x"00",  x"00",  x"00",  x"00",  x"b8",  x"9c",  x"a1",  x"9e", -- 1EA0
         x"9f",  x"00",  x"b5",  x"a7",  x"b3",  x"94",  x"a5",  x"a7", -- 1EA8
         x"6e",  x"a5",  x"ab",  x"00",  x"9e",  x"a7",  x"9e",  x"95", -- 1EB0
         x"9c",  x"50",  x"ba",  x"b5",  x"94",  x"00",  x"00",  x"00", -- 1EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED8
         x"00",  x"00",  x"00",  x"b8",  x"b3",  x"9d",  x"9e",  x"96", -- 1EE0
         x"94",  x"a5",  x"a1",  x"a4",  x"a2",  x"00",  x"b3",  x"b4", -- 1EE8
         x"ac",  x"a2",  x"a1",  x"00",  x"b7",  x"b5",  x"86",  x"9c", -- 1EF0
         x"50",  x"9c",  x"a4",  x"00",  x"6e",  x"00",  x"00",  x"00", -- 1EF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F38
         x"00",  x"00",  x"79",  x"78",  x"7b",  x"7a",  x"81",  x"78", -- 1F40
         x"93",  x"92",  x"91",  x"90",  x"8b",  x"8a",  x"7b",  x"7a", -- 1F48
         x"00",  x"88",  x"9a",  x"99",  x"79",  x"78",  x"83",  x"82", -- 1F50
         x"81",  x"78",  x"7b",  x"7a",  x"79",  x"78",  x"00",  x"00", -- 1F58
         x"00",  x"00",  x"75",  x"74",  x"77",  x"76",  x"7d",  x"7c", -- 1F60
         x"8f",  x"8e",  x"8d",  x"8c",  x"87",  x"84",  x"77",  x"76", -- 1F68
         x"85",  x"84",  x"98",  x"97",  x"75",  x"74",  x"7f",  x"7e", -- 1F70
         x"7d",  x"7c",  x"77",  x"76",  x"75",  x"74",  x"00",  x"00", -- 1F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
